��/  K��@AZ�����"SƤ`��g�o[j#ƽ�n-1��͈�P�Ǜ�*e�c�1��E#nT-�}����](0��'d���a�n�ƪ��H�.�1_�`1(WB>M�{*3��J�{|�S�&|}�@~H��c�9O�t�����}�n葥����29iY�IX����V�W|D&��1�^k��}��Tl�/*֍�����NX|���?�Q���`�C���q�43k�{tn�cVo $�$��q�W$�-��re �&{�s�B��>(y/nV���O���.s� �@J��Q�(��A@�C�q�*{������4��w�JL��y:���ҕ�@w�$�\��z��,��=0#�̑���0��Z��+�
��znY�+b��]Q���"�AX��s�3L̸e؉�9j�5�)��(=@NG���a�+R�q8�'R���^	d�$!���@�Q����Ww;M��VS� ��0Y�7%$i�,����>�lZ���PQ�[�Y�tɒ���r=����?�������p�g]�w���ên�q��JW�v�9K/b]����Q���Tt]@S�7�jx��� ��@@q�d�c��o&꯳��W��w�]H6���"�;�19�^v�A��$t����T�iǬ��P�>�[��1B��r��a=r��s#n9f�����*<Q�g`Sl�v��-��|�qtȉ%j���n�a��-ˑ�vMڏ��O�ѩu/c�\s2�E�)_D��/X��yg��-�/
��#@v�� ^��)�}间[��I�\D:3R9���J��Fg@*��oڂ׹L�H.�Q'L�����~�ϠX�/��n%{W�C�h]�A*a��	��;t~��\e-��5�ZJNND��� �0�%Ϗ
K���Hu�Dq0�Ā�����עD���B\����&�lW�vn���x�Ю�V�L�SV"��a5;^f�^�rV��h���Y<n�����@ay\��-ۯ�tؿ�)��l��.�45��1�gLl��B�M+G
�Y]���Bv�XU�=�[l������T��H
��=������8Ί
4��w7M2�N|���*�?�= YH��3��Ev��K����W�U���q�V����0y
�m�h��|g�i���CRS�o�]�M&?���L�G���68����U�G¡���~�y�In��>L8������`��M�#H��^D���A>g��dZ,���`;��q��5��>!w��4�
��-菴 ��ԥD1b㩴�6�r}+�9����x��eȻA�0���Bw��@9#3�ܹ���<S��9�\$����Ț��s�Ș�=`�)0��jD��� (��,�(�)̧�|�|P����zpǠ��\�i�M�&T���(�-9�g���P�w�Yv 7�](i|�?��G�b����|�W58�	]�lA��|2>Q2�j�˼"�&��@����� -n�Wd�U8�Z��F����H�.c�Ԧ�y��?�D ��5Wi�$���bB���6|/]B��r�.bu; װ�K����O�O��
�,��Y'��������c���V`r�L��W��N8bQ�\u��`1�.ռ�'��dE1:p��?�ڲ	N&�6S �ُ���Fas�U�hƙL�j֡a�C�3Dx���(���a�j@3_㉭mI&����F��E�g��DmrN�蝷k���\1����6%x��%O1���[9>����Y�e7t¤��!�=�A�Ҙ\.V�ة��هr���4���d��T,u�8����l�U�Nq�0�o�f����|��\ǐ�`�p�_(�v@���`cS8I�D���˪v��J�I��
����r����|��5���݅@���!bT���\co��S��a�/pt	lQ�77jU�I{k<)K�r#�����s#�1Ԕ�����_�֫��ْ�0��lxTYݜ�3f6r�0�Í7��d�D�t���vE٠g� Gk�<��~�i/����;�ئռ�a��8�G�f$ſP�ޗ�y���Ñ7V:	�����	^�\�O˴t��D�G;[FJH=�5J�R��v7�cB�p G�(����ܼmE�AТ�J�f_�+(ᛆ�!��v���iXA�\�RGfϡŀf�z�7��h�4��sd;5�`wA����j��RZT��#i+ �U�18�X�鄷_��������G|b����ϑd��{a@�*T1���&���2M��4�8
�5�V�#=�~d�(�U��.���^XBv:䡂Ѹ]�������쩫�:�.rx�E��V�N0l�a������7Dn��T�Mi����C�� u̩<]���/	(��Q����������w����fj����*8b��0���j�Ie��A����'��|"ɕ��{���� {w��6e�v򆒯��h��Y�g�fe�C���8
�K}S俿G��C�rꮩ�z�D}�)tO���/��5}Ă>h�OgA�	]��LZc��)O���ʌNz��+4|�G4c+�f�N>� [�����ǲ�샲��!���hF|h8�|�;��!��7c�j�4�����<��p�s�6��ݠsX�τlhǯ�&����^���O}S���$ڨ�Kk�����M��;�7ȳ�Y[��lU-�(r��Z��WstJO��3��_=��zq=r}64w^΄��:����s�b�K��; ̇�&(
�1R�sQ�9AWݰ��;�9K�����yR$�;��T�S�2l9��h^�^��x@T*Ba`iP�Iۯ�]��y��.�S��ŕ��V:�@+�C��|��;={w8`���B�~�ik��p��/M�4r"��P���hr/
�['oj`�$}I�We���^�}����&*��1� �ᎴK�xSP��E8BX��/�7��x/���&ـ8�g��q��ѿ2 ����۩�R��@�iy%~l�.�r�t�7�̓ rs���̎v�j�Y�jT�@�a"ߢZ�E91����̢��X����i�Ì��\!Z�h�Rr��+��{K�w�u�,�L���t�g��a�Y@��Z1� �����i�(��l,�	�l��߿���Z�B��R��������'Y���H����$�dz�1�Xu���~��3�o�K��\H�x
6V�-�@���D��~�p��j�*��]8!^�hccX��m6�I>-�� �LY�U��3 ��#�h��f	wO!�� 8�������C��{�\���񾧯�#P��+u�!�'۽w�2���и��Q�a�A$��>|Rl�ps�,�&��J�(z(ɥ��ҩ�5ȏY�A?,s�&����J�,�	�� �z���ӈ,aez�0�"��S`�a��Hm�db����ֶD˻ʠف�;�C�M�4q�=&ޭ�f��5�h��{����J)
��c�*VpG��.wY�f���U'�ЮÒ��̑��4��?*���������C��V[u� ���������=r�y�^l@s7v1��s