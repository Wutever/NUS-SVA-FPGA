// de2_115_WEB_Qsys.v

// Generated using ACDS version 12.0 178 at 2017.06.29.23:56:58

`timescale 1 ps / 1 ps
module de2_115_WEB_Qsys (
		output wire        sd_clk_external_connection_export,                               //          sd_clk_external_connection.export
		inout  wire        i2c_sda_external_connection_export,                              //         i2c_sda_external_connection.export
		output wire        altpll_c1_clk,                                                   //                           altpll_c1.clk
		inout  wire [3:0]  sd_dat_external_connection_export,                               //          sd_dat_external_connection.export
		inout  wire [7:0]  lcd_external_data,                                               //                        lcd_external.data
		output wire        lcd_external_E,                                                  //                                    .E
		output wire        lcd_external_RS,                                                 //                                    .RS
		output wire        lcd_external_RW,                                                 //                                    .RW
		output wire        altpll_c3_clk,                                                   //                           altpll_c3.clk
		output wire        c2_out_clk_clk,                                                  //                          c2_out_clk.clk
		inout  wire        epp_i2c_sda_external_connection_export,                          //     epp_i2c_sda_external_connection.export
		output wire        altpll_phasedone_conduit_export,                                 //            altpll_phasedone_conduit.export
		output wire        i2c_scl_external_connection_export,                              //         i2c_scl_external_connection.export
		output wire [8:0]  ledg_external_connection_export,                                 //            ledg_external_connection.export
		output wire        c0_out_clk_clk,                                                  //                          c0_out_clk.clk
		output wire        audio_conduit_end_XCK,                                           //                   audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,                                        //                                    .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,                                        //                                    .ADCLRC
		output wire        audio_conduit_end_DACDAT,                                        //                                    .DACDAT
		input  wire        audio_conduit_end_DACLRC,                                        //                                    .DACLRC
		input  wire        audio_conduit_end_BCLK,                                          //                                    .BCLK
		input  wire        reset_reset_n,                                                   //                               reset.reset_n
		output wire [22:0] tri_state_bridge_flash_bridge_0_out_address_to_the_cfi_flash,    // tri_state_bridge_flash_bridge_0_out.address_to_the_cfi_flash
		inout  wire [7:0]  tri_state_bridge_flash_bridge_0_out_tri_state_bridge_flash_data, //                                    .tri_state_bridge_flash_data
		output wire [0:0]  tri_state_bridge_flash_bridge_0_out_write_n_to_the_cfi_flash,    //                                    .write_n_to_the_cfi_flash
		output wire [0:0]  tri_state_bridge_flash_bridge_0_out_select_n_to_the_cfi_flash,   //                                    .select_n_to_the_cfi_flash
		output wire [0:0]  tri_state_bridge_flash_bridge_0_out_read_n_to_the_cfi_flash,     //                                    .read_n_to_the_cfi_flash
		input  wire        rs232_external_connection_rxd,                                   //           rs232_external_connection.rxd
		output wire        rs232_external_connection_txd,                                   //                                    .txd
		input  wire        rs232_external_connection_cts_n,                                 //                                    .cts_n
		output wire        rs232_external_connection_rts_n,                                 //                                    .rts_n
		input  wire        ir_external_connection_export,                                   //              ir_external_connection.export
		input  wire [3:0]  tse_mac_conduit_connection_m_rx_d,                               //          tse_mac_conduit_connection.m_rx_d
		input  wire        tse_mac_conduit_connection_m_rx_en,                              //                                    .m_rx_en
		input  wire        tse_mac_conduit_connection_m_rx_err,                             //                                    .m_rx_err
		output wire [3:0]  tse_mac_conduit_connection_m_tx_d,                               //                                    .m_tx_d
		output wire        tse_mac_conduit_connection_m_tx_en,                              //                                    .m_tx_en
		output wire        tse_mac_conduit_connection_m_tx_err,                             //                                    .m_tx_err
		input  wire        tse_mac_conduit_connection_tx_clk,                               //                                    .tx_clk
		input  wire        tse_mac_conduit_connection_rx_clk,                               //                                    .rx_clk
		input  wire        tse_mac_conduit_connection_set_10,                               //                                    .set_10
		input  wire        tse_mac_conduit_connection_set_1000,                             //                                    .set_1000
		output wire        tse_mac_conduit_connection_ena_10,                               //                                    .ena_10
		output wire        tse_mac_conduit_connection_eth_mode,                             //                                    .eth_mode
		output wire        tse_mac_conduit_connection_mdio_out,                             //                                    .mdio_out
		output wire        tse_mac_conduit_connection_mdio_oen,                             //                                    .mdio_oen
		input  wire        tse_mac_conduit_connection_mdio_in,                              //                                    .mdio_in
		output wire        tse_mac_conduit_connection_mdc,                                  //                                    .mdc
		input  wire        tse_mac_conduit_connection_m_rx_col,                             //                                    .m_rx_col
		input  wire        tse_mac_conduit_connection_m_rx_crs,                             //                                    .m_rx_crs
		output wire        sma_out_external_connection_export,                              //         sma_out_external_connection.export
		input  wire [3:0]  key_external_connection_export,                                  //             key_external_connection.export
		inout  wire [15:0] isp1362_if_0_conduit_end_DATA,                                   //            isp1362_if_0_conduit_end.DATA
		output wire [1:0]  isp1362_if_0_conduit_end_ADDR,                                   //                                    .ADDR
		output wire        isp1362_if_0_conduit_end_RD_N,                                   //                                    .RD_N
		output wire        isp1362_if_0_conduit_end_WR_N,                                   //                                    .WR_N
		output wire        isp1362_if_0_conduit_end_CS_N,                                   //                                    .CS_N
		output wire        isp1362_if_0_conduit_end_RST_N,                                  //                                    .RST_N
		input  wire        isp1362_if_0_conduit_end_INT0,                                   //                                    .INT0
		input  wire        isp1362_if_0_conduit_end_INT1,                                   //                                    .INT1
		input  wire        clk_50_clk_in_clk,                                               //                       clk_50_clk_in.clk
		output wire        altpll_locked_conduit_export,                                    //               altpll_locked_conduit.export
		output wire        epp_i2c_scl_external_connection_export,                          //     epp_i2c_scl_external_connection.export
		inout  wire [15:0] sram_conduit_end_DQ,                                             //                    sram_conduit_end.DQ
		output wire [19:0] sram_conduit_end_ADDR,                                           //                                    .ADDR
		output wire        sram_conduit_end_UB_n,                                           //                                    .UB_n
		output wire        sram_conduit_end_LB_n,                                           //                                    .LB_n
		output wire        sram_conduit_end_WE_n,                                           //                                    .WE_n
		output wire        sram_conduit_end_CE_n,                                           //                                    .CE_n
		output wire        sram_conduit_end_OE_n,                                           //                                    .OE_n
		input  wire        sd_wp_n_external_connection_export,                              //         sd_wp_n_external_connection.export
		input  wire        sma_in_external_connection_export,                               //          sma_in_external_connection.export
		input  wire        clkoutput_export,                                                //                           clkoutput.export
		input  wire        altpll_areset_conduit_export,                                    //               altpll_areset_conduit.export
		output wire [63:0] seg7_conduit_end_export,                                         //                    seg7_conduit_end.export
		output wire [12:0] sdram_wire_addr,                                                 //                          sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                                   //                                    .ba
		output wire        sdram_wire_cas_n,                                                //                                    .cas_n
		output wire        sdram_wire_cke,                                                  //                                    .cke
		output wire        sdram_wire_cs_n,                                                 //                                    .cs_n
		inout  wire [31:0] sdram_wire_dq,                                                   //                                    .dq
		output wire [3:0]  sdram_wire_dqm,                                                  //                                    .dqm
		output wire        sdram_wire_ras_n,                                                //                                    .ras_n
		output wire        sdram_wire_we_n,                                                 //                                    .we_n
		input  wire [13:0] dataoutput_export,                                               //                          dataoutput.export
		input  wire [17:0] sw_external_connection_export,                                   //              sw_external_connection.export
		output wire [17:0] ledr_external_connection_export,                                 //            ledr_external_connection.export
		inout  wire        sd_cmd_external_connection_export                                //          sd_cmd_external_connection.export
	);

	wire    [7:0] tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in;                            // tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_in -> tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data_in
	wire    [7:0] tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out;                           // tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data
	wire          tri_state_flash_bridge_pinsharer_0_tcm_grant;                                                     // tri_state_bridge_flash_bridge_0:grant -> tri_state_flash_bridge_pinSharer_0:grant
	wire    [0:0] tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out;                             // tri_state_flash_bridge_pinSharer_0:select_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_select_n_to_the_cfi_flash
	wire          tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen;                         // tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data_outen -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_outen
	wire          tri_state_flash_bridge_pinsharer_0_tcm_request;                                                   // tri_state_flash_bridge_pinSharer_0:request -> tri_state_bridge_flash_bridge_0:request
	wire    [0:0] tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out;                              // tri_state_flash_bridge_pinSharer_0:write_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_write_n_to_the_cfi_flash
	wire    [0:0] tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out;                               // tri_state_flash_bridge_pinSharer_0:read_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_read_n_to_the_cfi_flash
	wire   [22:0] tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out;                              // tri_state_flash_bridge_pinSharer_0:address_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_address_to_the_cfi_flash
	wire          cfi_flash_tcm_chipselect_n_out;                                                                   // cfi_flash:tcm_chipselect_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_chipselect_n_out
	wire          cfi_flash_tcm_grant;                                                                              // tri_state_flash_bridge_pinSharer_0:tcs0_grant -> cfi_flash:tcm_grant
	wire          cfi_flash_tcm_data_outen;                                                                         // cfi_flash:tcm_data_outen -> tri_state_flash_bridge_pinSharer_0:tcs0_data_outen
	wire          cfi_flash_tcm_request;                                                                            // cfi_flash:tcm_request -> tri_state_flash_bridge_pinSharer_0:tcs0_request
	wire    [7:0] cfi_flash_tcm_data_out;                                                                           // cfi_flash:tcm_data_out -> tri_state_flash_bridge_pinSharer_0:tcs0_data_out
	wire          cfi_flash_tcm_write_n_out;                                                                        // cfi_flash:tcm_write_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_write_n_out
	wire   [22:0] cfi_flash_tcm_address_out;                                                                        // cfi_flash:tcm_address_out -> tri_state_flash_bridge_pinSharer_0:tcs0_address_out
	wire    [7:0] cfi_flash_tcm_data_in;                                                                            // tri_state_flash_bridge_pinSharer_0:tcs0_data_in -> cfi_flash:tcm_data_in
	wire          cfi_flash_tcm_read_n_out;                                                                         // cfi_flash:tcm_read_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_read_n_out
	wire          cpu_jtag_debug_module_reset_reset;                                                                // cpu:jtag_debug_module_resetrequest -> [ISP1362_IF_0:avs_dc_reset_n_iRST_N, ISP1362_IF_0_dc_translator:reset, ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:reset, ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_011:reset, rsp_xbar_demux_011:reset, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	wire          tse_mac_receive_endofpacket;                                                                      // tse_mac:ff_rx_eop -> sgdma_rx:in_endofpacket
	wire          tse_mac_receive_valid;                                                                            // tse_mac:ff_rx_dval -> sgdma_rx:in_valid
	wire          tse_mac_receive_startofpacket;                                                                    // tse_mac:ff_rx_sop -> sgdma_rx:in_startofpacket
	wire    [5:0] tse_mac_receive_error;                                                                            // tse_mac:rx_err -> sgdma_rx:in_error
	wire    [1:0] tse_mac_receive_empty;                                                                            // tse_mac:ff_rx_mod -> sgdma_rx:in_empty
	wire   [31:0] tse_mac_receive_data;                                                                             // tse_mac:ff_rx_data -> sgdma_rx:in_data
	wire          tse_mac_receive_ready;                                                                            // sgdma_rx:in_ready -> tse_mac:ff_rx_rdy
	wire          sgdma_tx_out_endofpacket;                                                                         // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire          sgdma_tx_out_valid;                                                                               // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire          sgdma_tx_out_startofpacket;                                                                       // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire          sgdma_tx_out_error;                                                                               // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire    [1:0] sgdma_tx_out_empty;                                                                               // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire   [31:0] sgdma_tx_out_data;                                                                                // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire          sgdma_tx_out_ready;                                                                               // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire          cpu_instruction_master_waitrequest;                                                               // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [27:0] cpu_instruction_master_address;                                                                   // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                      // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                  // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                             // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire          cpu_data_master_waitrequest;                                                                      // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                        // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [27:0] cpu_data_master_address;                                                                          // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                            // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                             // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                         // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                      // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire          cpu_data_master_readdatavalid;                                                                    // cpu_data_master_translator:av_readdatavalid -> cpu:d_readdatavalid
	wire    [3:0] cpu_data_master_byteenable;                                                                       // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          sgdma_tx_descriptor_read_waitrequest;                                                             // sgdma_tx_descriptor_read_translator:av_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire   [31:0] sgdma_tx_descriptor_read_address;                                                                 // sgdma_tx:descriptor_read_address -> sgdma_tx_descriptor_read_translator:av_address
	wire          sgdma_tx_descriptor_read_read;                                                                    // sgdma_tx:descriptor_read_read -> sgdma_tx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_tx_descriptor_read_readdata;                                                                // sgdma_tx_descriptor_read_translator:av_readdata -> sgdma_tx:descriptor_read_readdata
	wire          sgdma_tx_descriptor_read_readdatavalid;                                                           // sgdma_tx_descriptor_read_translator:av_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire          sgdma_tx_descriptor_write_waitrequest;                                                            // sgdma_tx_descriptor_write_translator:av_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire   [31:0] sgdma_tx_descriptor_write_writedata;                                                              // sgdma_tx:descriptor_write_writedata -> sgdma_tx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_address;                                                                // sgdma_tx:descriptor_write_address -> sgdma_tx_descriptor_write_translator:av_address
	wire          sgdma_tx_descriptor_write_write;                                                                  // sgdma_tx:descriptor_write_write -> sgdma_tx_descriptor_write_translator:av_write
	wire          sgdma_rx_descriptor_read_waitrequest;                                                             // sgdma_rx_descriptor_read_translator:av_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire   [31:0] sgdma_rx_descriptor_read_address;                                                                 // sgdma_rx:descriptor_read_address -> sgdma_rx_descriptor_read_translator:av_address
	wire          sgdma_rx_descriptor_read_read;                                                                    // sgdma_rx:descriptor_read_read -> sgdma_rx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_rx_descriptor_read_readdata;                                                                // sgdma_rx_descriptor_read_translator:av_readdata -> sgdma_rx:descriptor_read_readdata
	wire          sgdma_rx_descriptor_read_readdatavalid;                                                           // sgdma_rx_descriptor_read_translator:av_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire          sgdma_rx_descriptor_write_waitrequest;                                                            // sgdma_rx_descriptor_write_translator:av_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire   [31:0] sgdma_rx_descriptor_write_writedata;                                                              // sgdma_rx:descriptor_write_writedata -> sgdma_rx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_address;                                                                // sgdma_rx:descriptor_write_address -> sgdma_rx_descriptor_write_translator:av_address
	wire          sgdma_rx_descriptor_write_write;                                                                  // sgdma_rx:descriptor_write_write -> sgdma_rx_descriptor_write_translator:av_write
	wire          sgdma_tx_m_read_waitrequest;                                                                      // sgdma_tx_m_read_translator:av_waitrequest -> sgdma_tx:m_read_waitrequest
	wire   [31:0] sgdma_tx_m_read_address;                                                                          // sgdma_tx:m_read_address -> sgdma_tx_m_read_translator:av_address
	wire          sgdma_tx_m_read_read;                                                                             // sgdma_tx:m_read_read -> sgdma_tx_m_read_translator:av_read
	wire   [31:0] sgdma_tx_m_read_readdata;                                                                         // sgdma_tx_m_read_translator:av_readdata -> sgdma_tx:m_read_readdata
	wire          sgdma_tx_m_read_readdatavalid;                                                                    // sgdma_tx_m_read_translator:av_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire          sgdma_rx_m_write_waitrequest;                                                                     // sgdma_rx_m_write_translator:av_waitrequest -> sgdma_rx:m_write_waitrequest
	wire   [31:0] sgdma_rx_m_write_writedata;                                                                       // sgdma_rx:m_write_writedata -> sgdma_rx_m_write_translator:av_writedata
	wire   [31:0] sgdma_rx_m_write_address;                                                                         // sgdma_rx:m_write_address -> sgdma_rx_m_write_translator:av_address
	wire          sgdma_rx_m_write_write;                                                                           // sgdma_rx:m_write_write -> sgdma_rx_m_write_translator:av_write
	wire    [3:0] sgdma_rx_m_write_byteenable;                                                                      // sgdma_rx:m_write_byteenable -> sgdma_rx_m_write_translator:av_byteenable
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_jtag_debug_module_translator:av_chipselect -> cpu:jtag_debug_module_select
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_jtag_debug_module_translator:av_begintransfer -> cpu:jtag_debug_module_begintransfer
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_waitrequest;                                         // cfi_flash:uas_waitrequest -> cfi_flash_uas_translator:av_waitrequest
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_burstcount;                                          // cfi_flash_uas_translator:av_burstcount -> cfi_flash:uas_burstcount
	wire    [7:0] cfi_flash_uas_translator_avalon_anti_slave_0_writedata;                                           // cfi_flash_uas_translator:av_writedata -> cfi_flash:uas_writedata
	wire   [22:0] cfi_flash_uas_translator_avalon_anti_slave_0_address;                                             // cfi_flash_uas_translator:av_address -> cfi_flash:uas_address
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_lock;                                                // cfi_flash_uas_translator:av_lock -> cfi_flash:uas_lock
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_write;                                               // cfi_flash_uas_translator:av_write -> cfi_flash:uas_write
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_read;                                                // cfi_flash_uas_translator:av_read -> cfi_flash:uas_read
	wire    [7:0] cfi_flash_uas_translator_avalon_anti_slave_0_readdata;                                            // cfi_flash:uas_readdata -> cfi_flash_uas_translator:av_readdata
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_debugaccess;                                         // cfi_flash_uas_translator:av_debugaccess -> cfi_flash:uas_debugaccess
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_readdatavalid;                                       // cfi_flash:uas_readdatavalid -> cfi_flash_uas_translator:av_readdatavalid
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_byteenable;                                          // cfi_flash_uas_translator:av_byteenable -> cfi_flash:uas_byteenable
	wire   [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_writedata;                                       // onchip_memory2_s1_translator:av_writedata -> onchip_memory2:writedata
	wire   [14:0] onchip_memory2_s1_translator_avalon_anti_slave_0_address;                                         // onchip_memory2_s1_translator:av_address -> onchip_memory2:address
	wire          onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect;                                      // onchip_memory2_s1_translator:av_chipselect -> onchip_memory2:chipselect
	wire          onchip_memory2_s1_translator_avalon_anti_slave_0_clken;                                           // onchip_memory2_s1_translator:av_clken -> onchip_memory2:clken
	wire          onchip_memory2_s1_translator_avalon_anti_slave_0_write;                                           // onchip_memory2_s1_translator:av_write -> onchip_memory2:write
	wire   [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_readdata;                                        // onchip_memory2:readdata -> onchip_memory2_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable;                                      // onchip_memory2_s1_translator:av_byteenable -> onchip_memory2:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                              // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [24:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                  // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                               // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                    // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                     // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                 // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                            // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [3:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                               // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [15:0] sram_avalon_slave_translator_avalon_anti_slave_0_writedata;                                       // sram_avalon_slave_translator:av_writedata -> sram:s_writedata
	wire   [19:0] sram_avalon_slave_translator_avalon_anti_slave_0_address;                                         // sram_avalon_slave_translator:av_address -> sram:s_address
	wire          sram_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                      // sram_avalon_slave_translator:av_chipselect -> sram:s_chipselect_n
	wire          sram_avalon_slave_translator_avalon_anti_slave_0_write;                                           // sram_avalon_slave_translator:av_write -> sram:s_write_n
	wire          sram_avalon_slave_translator_avalon_anti_slave_0_read;                                            // sram_avalon_slave_translator:av_read -> sram:s_read_n
	wire   [15:0] sram_avalon_slave_translator_avalon_anti_slave_0_readdata;                                        // sram:s_readdata -> sram_avalon_slave_translator:av_readdata
	wire    [1:0] sram_avalon_slave_translator_avalon_anti_slave_0_byteenable;                                      // sram_avalon_slave_translator:av_byteenable -> sram:s_byteenable_n
	wire          clock_crossing_io_s0_translator_avalon_anti_slave_0_waitrequest;                                  // clock_crossing_io:s0_waitrequest -> clock_crossing_io_s0_translator:av_waitrequest
	wire          clock_crossing_io_s0_translator_avalon_anti_slave_0_burstcount;                                   // clock_crossing_io_s0_translator:av_burstcount -> clock_crossing_io:s0_burstcount
	wire   [31:0] clock_crossing_io_s0_translator_avalon_anti_slave_0_writedata;                                    // clock_crossing_io_s0_translator:av_writedata -> clock_crossing_io:s0_writedata
	wire    [8:0] clock_crossing_io_s0_translator_avalon_anti_slave_0_address;                                      // clock_crossing_io_s0_translator:av_address -> clock_crossing_io:s0_address
	wire          clock_crossing_io_s0_translator_avalon_anti_slave_0_write;                                        // clock_crossing_io_s0_translator:av_write -> clock_crossing_io:s0_write
	wire          clock_crossing_io_s0_translator_avalon_anti_slave_0_read;                                         // clock_crossing_io_s0_translator:av_read -> clock_crossing_io:s0_read
	wire   [31:0] clock_crossing_io_s0_translator_avalon_anti_slave_0_readdata;                                     // clock_crossing_io:s0_readdata -> clock_crossing_io_s0_translator:av_readdata
	wire          clock_crossing_io_s0_translator_avalon_anti_slave_0_debugaccess;                                  // clock_crossing_io_s0_translator:av_debugaccess -> clock_crossing_io:s0_debugaccess
	wire          clock_crossing_io_s0_translator_avalon_anti_slave_0_readdatavalid;                                // clock_crossing_io:s0_readdatavalid -> clock_crossing_io_s0_translator:av_readdatavalid
	wire    [3:0] clock_crossing_io_s0_translator_avalon_anti_slave_0_byteenable;                                   // clock_crossing_io_s0_translator:av_byteenable -> clock_crossing_io:s0_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] audio_avalon_slave_translator_avalon_anti_slave_0_writedata;                                      // audio_avalon_slave_translator:av_writedata -> audio:avs_s1_writedata
	wire    [2:0] audio_avalon_slave_translator_avalon_anti_slave_0_address;                                        // audio_avalon_slave_translator:av_address -> audio:avs_s1_address
	wire          audio_avalon_slave_translator_avalon_anti_slave_0_write;                                          // audio_avalon_slave_translator:av_write -> audio:avs_s1_write
	wire          audio_avalon_slave_translator_avalon_anti_slave_0_read;                                           // audio_avalon_slave_translator:av_read -> audio:avs_s1_read
	wire   [15:0] audio_avalon_slave_translator_avalon_anti_slave_0_readdata;                                       // audio:avs_s1_readdata -> audio_avalon_slave_translator:av_readdata
	wire   [31:0] altpll_pll_slave_translator_avalon_anti_slave_0_writedata;                                        // altpll_pll_slave_translator:av_writedata -> altpll:writedata
	wire    [1:0] altpll_pll_slave_translator_avalon_anti_slave_0_address;                                          // altpll_pll_slave_translator:av_address -> altpll:address
	wire          altpll_pll_slave_translator_avalon_anti_slave_0_write;                                            // altpll_pll_slave_translator:av_write -> altpll:write
	wire          altpll_pll_slave_translator_avalon_anti_slave_0_read;                                             // altpll_pll_slave_translator:av_read -> altpll:read
	wire   [31:0] altpll_pll_slave_translator_avalon_anti_slave_0_readdata;                                         // altpll:readdata -> altpll_pll_slave_translator:av_readdata
	wire    [1:0] sma_in_s1_translator_avalon_anti_slave_0_address;                                                 // sma_in_s1_translator:av_address -> sma_in:address
	wire   [31:0] sma_in_s1_translator_avalon_anti_slave_0_readdata;                                                // sma_in:readdata -> sma_in_s1_translator:av_readdata
	wire   [31:0] sma_out_s1_translator_avalon_anti_slave_0_writedata;                                              // sma_out_s1_translator:av_writedata -> sma_out:writedata
	wire    [1:0] sma_out_s1_translator_avalon_anti_slave_0_address;                                                // sma_out_s1_translator:av_address -> sma_out:address
	wire          sma_out_s1_translator_avalon_anti_slave_0_chipselect;                                             // sma_out_s1_translator:av_chipselect -> sma_out:chipselect
	wire          sma_out_s1_translator_avalon_anti_slave_0_write;                                                  // sma_out_s1_translator:av_write -> sma_out:write_n
	wire   [31:0] sma_out_s1_translator_avalon_anti_slave_0_readdata;                                               // sma_out:readdata -> sma_out_s1_translator:av_readdata
	wire   [15:0] isp1362_if_0_dc_translator_avalon_anti_slave_0_writedata;                                         // ISP1362_IF_0_dc_translator:av_writedata -> ISP1362_IF_0:avs_dc_writedata_iDATA
	wire          isp1362_if_0_dc_translator_avalon_anti_slave_0_address;                                           // ISP1362_IF_0_dc_translator:av_address -> ISP1362_IF_0:avs_dc_address_iADDR
	wire          isp1362_if_0_dc_translator_avalon_anti_slave_0_chipselect;                                        // ISP1362_IF_0_dc_translator:av_chipselect -> ISP1362_IF_0:avs_dc_chipselect_n_iCS_N
	wire          isp1362_if_0_dc_translator_avalon_anti_slave_0_write;                                             // ISP1362_IF_0_dc_translator:av_write -> ISP1362_IF_0:avs_dc_write_n_iWR_N
	wire          isp1362_if_0_dc_translator_avalon_anti_slave_0_read;                                              // ISP1362_IF_0_dc_translator:av_read -> ISP1362_IF_0:avs_dc_read_n_iRD_N
	wire   [15:0] isp1362_if_0_dc_translator_avalon_anti_slave_0_readdata;                                          // ISP1362_IF_0:avs_dc_readdata_oDATA -> ISP1362_IF_0_dc_translator:av_readdata
	wire   [15:0] isp1362_if_0_hc_translator_avalon_anti_slave_0_writedata;                                         // ISP1362_IF_0_hc_translator:av_writedata -> ISP1362_IF_0:avs_hc_writedata_iDATA
	wire          isp1362_if_0_hc_translator_avalon_anti_slave_0_address;                                           // ISP1362_IF_0_hc_translator:av_address -> ISP1362_IF_0:avs_hc_address_iADDR
	wire          isp1362_if_0_hc_translator_avalon_anti_slave_0_chipselect;                                        // ISP1362_IF_0_hc_translator:av_chipselect -> ISP1362_IF_0:avs_hc_chipselect_n_iCS_N
	wire          isp1362_if_0_hc_translator_avalon_anti_slave_0_write;                                             // ISP1362_IF_0_hc_translator:av_write -> ISP1362_IF_0:avs_hc_write_n_iWR_N
	wire          isp1362_if_0_hc_translator_avalon_anti_slave_0_read;                                              // ISP1362_IF_0_hc_translator:av_read -> ISP1362_IF_0:avs_hc_read_n_iRD_N
	wire   [15:0] isp1362_if_0_hc_translator_avalon_anti_slave_0_readdata;                                          // ISP1362_IF_0:avs_hc_readdata_oDATA -> ISP1362_IF_0_hc_translator:av_readdata
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_writedata;                                    // descriptor_memory_s1_translator:av_writedata -> descriptor_memory:writedata
	wire    [9:0] descriptor_memory_s1_translator_avalon_anti_slave_0_address;                                      // descriptor_memory_s1_translator:av_address -> descriptor_memory:address
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect;                                   // descriptor_memory_s1_translator:av_chipselect -> descriptor_memory:chipselect
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_clken;                                        // descriptor_memory_s1_translator:av_clken -> descriptor_memory:clken
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_write;                                        // descriptor_memory_s1_translator:av_write -> descriptor_memory:write
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_readdata;                                     // descriptor_memory:readdata -> descriptor_memory_s1_translator:av_readdata
	wire    [3:0] descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable;                                   // descriptor_memory_s1_translator:av_byteenable -> descriptor_memory:byteenable
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_writedata;                                            // sgdma_rx_csr_translator:av_writedata -> sgdma_rx:csr_writedata
	wire    [3:0] sgdma_rx_csr_translator_avalon_anti_slave_0_address;                                              // sgdma_rx_csr_translator:av_address -> sgdma_rx:csr_address
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect;                                           // sgdma_rx_csr_translator:av_chipselect -> sgdma_rx:csr_chipselect
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_write;                                                // sgdma_rx_csr_translator:av_write -> sgdma_rx:csr_write
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_read;                                                 // sgdma_rx_csr_translator:av_read -> sgdma_rx:csr_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_readdata;                                             // sgdma_rx:csr_readdata -> sgdma_rx_csr_translator:av_readdata
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_writedata;                                            // sgdma_tx_csr_translator:av_writedata -> sgdma_tx:csr_writedata
	wire    [3:0] sgdma_tx_csr_translator_avalon_anti_slave_0_address;                                              // sgdma_tx_csr_translator:av_address -> sgdma_tx:csr_address
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect;                                           // sgdma_tx_csr_translator:av_chipselect -> sgdma_tx:csr_chipselect
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_write;                                                // sgdma_tx_csr_translator:av_write -> sgdma_tx:csr_write
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_read;                                                 // sgdma_tx_csr_translator:av_read -> sgdma_tx:csr_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_readdata;                                             // sgdma_tx:csr_readdata -> sgdma_tx_csr_translator:av_readdata
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest;                                  // tse_mac:waitrequest -> tse_mac_control_port_translator:av_waitrequest
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_writedata;                                    // tse_mac_control_port_translator:av_writedata -> tse_mac:writedata
	wire    [7:0] tse_mac_control_port_translator_avalon_anti_slave_0_address;                                      // tse_mac_control_port_translator:av_address -> tse_mac:address
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_write;                                        // tse_mac_control_port_translator:av_write -> tse_mac:write
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_read;                                         // tse_mac_control_port_translator:av_read -> tse_mac:read
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_readdata;                                     // tse_mac:readdata -> tse_mac_control_port_translator:av_readdata
	wire    [1:0] pio_0_s1_translator_avalon_anti_slave_0_address;                                                  // pio_0_s1_translator:av_address -> pio_0:address
	wire   [31:0] pio_0_s1_translator_avalon_anti_slave_0_readdata;                                                 // pio_0:readdata -> pio_0_s1_translator:av_readdata
	wire    [1:0] pio_1_s1_translator_avalon_anti_slave_0_address;                                                  // pio_1_s1_translator:av_address -> pio_1:address
	wire   [31:0] pio_1_s1_translator_avalon_anti_slave_0_readdata;                                                 // pio_1:readdata -> pio_1_s1_translator:av_readdata
	wire    [0:0] clock_crossing_io_m0_burstcount;                                                                  // clock_crossing_io:m0_burstcount -> clock_crossing_io_m0_translator:av_burstcount
	wire          clock_crossing_io_m0_waitrequest;                                                                 // clock_crossing_io_m0_translator:av_waitrequest -> clock_crossing_io:m0_waitrequest
	wire    [8:0] clock_crossing_io_m0_address;                                                                     // clock_crossing_io:m0_address -> clock_crossing_io_m0_translator:av_address
	wire   [31:0] clock_crossing_io_m0_writedata;                                                                   // clock_crossing_io:m0_writedata -> clock_crossing_io_m0_translator:av_writedata
	wire          clock_crossing_io_m0_write;                                                                       // clock_crossing_io:m0_write -> clock_crossing_io_m0_translator:av_write
	wire          clock_crossing_io_m0_read;                                                                        // clock_crossing_io:m0_read -> clock_crossing_io_m0_translator:av_read
	wire   [31:0] clock_crossing_io_m0_readdata;                                                                    // clock_crossing_io_m0_translator:av_readdata -> clock_crossing_io:m0_readdata
	wire          clock_crossing_io_m0_debugaccess;                                                                 // clock_crossing_io:m0_debugaccess -> clock_crossing_io_m0_translator:av_debugaccess
	wire    [3:0] clock_crossing_io_m0_byteenable;                                                                  // clock_crossing_io:m0_byteenable -> clock_crossing_io_m0_translator:av_byteenable
	wire          clock_crossing_io_m0_readdatavalid;                                                               // clock_crossing_io_m0_translator:av_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire   [31:0] key_s1_translator_avalon_anti_slave_0_writedata;                                                  // key_s1_translator:av_writedata -> key:writedata
	wire    [1:0] key_s1_translator_avalon_anti_slave_0_address;                                                    // key_s1_translator:av_address -> key:address
	wire          key_s1_translator_avalon_anti_slave_0_chipselect;                                                 // key_s1_translator:av_chipselect -> key:chipselect
	wire          key_s1_translator_avalon_anti_slave_0_write;                                                      // key_s1_translator:av_write -> key:write_n
	wire   [31:0] key_s1_translator_avalon_anti_slave_0_readdata;                                                   // key:readdata -> key_s1_translator:av_readdata
	wire    [7:0] lcd_control_slave_translator_avalon_anti_slave_0_writedata;                                       // lcd_control_slave_translator:av_writedata -> lcd:writedata
	wire    [1:0] lcd_control_slave_translator_avalon_anti_slave_0_address;                                         // lcd_control_slave_translator:av_address -> lcd:address
	wire          lcd_control_slave_translator_avalon_anti_slave_0_write;                                           // lcd_control_slave_translator:av_write -> lcd:write
	wire          lcd_control_slave_translator_avalon_anti_slave_0_read;                                            // lcd_control_slave_translator:av_read -> lcd:read
	wire    [7:0] lcd_control_slave_translator_avalon_anti_slave_0_readdata;                                        // lcd:readdata -> lcd_control_slave_translator:av_readdata
	wire          lcd_control_slave_translator_avalon_anti_slave_0_begintransfer;                                   // lcd_control_slave_translator:av_begintransfer -> lcd:begintransfer
	wire   [31:0] sd_clk_s1_translator_avalon_anti_slave_0_writedata;                                               // sd_clk_s1_translator:av_writedata -> sd_clk:writedata
	wire    [1:0] sd_clk_s1_translator_avalon_anti_slave_0_address;                                                 // sd_clk_s1_translator:av_address -> sd_clk:address
	wire          sd_clk_s1_translator_avalon_anti_slave_0_chipselect;                                              // sd_clk_s1_translator:av_chipselect -> sd_clk:chipselect
	wire          sd_clk_s1_translator_avalon_anti_slave_0_write;                                                   // sd_clk_s1_translator:av_write -> sd_clk:write_n
	wire   [31:0] sd_clk_s1_translator_avalon_anti_slave_0_readdata;                                                // sd_clk:readdata -> sd_clk_s1_translator:av_readdata
	wire   [31:0] sd_cmd_s1_translator_avalon_anti_slave_0_writedata;                                               // sd_cmd_s1_translator:av_writedata -> sd_cmd:writedata
	wire    [1:0] sd_cmd_s1_translator_avalon_anti_slave_0_address;                                                 // sd_cmd_s1_translator:av_address -> sd_cmd:address
	wire          sd_cmd_s1_translator_avalon_anti_slave_0_chipselect;                                              // sd_cmd_s1_translator:av_chipselect -> sd_cmd:chipselect
	wire          sd_cmd_s1_translator_avalon_anti_slave_0_write;                                                   // sd_cmd_s1_translator:av_write -> sd_cmd:write_n
	wire   [31:0] sd_cmd_s1_translator_avalon_anti_slave_0_readdata;                                                // sd_cmd:readdata -> sd_cmd_s1_translator:av_readdata
	wire   [31:0] sd_dat_s1_translator_avalon_anti_slave_0_writedata;                                               // sd_dat_s1_translator:av_writedata -> sd_dat:writedata
	wire    [1:0] sd_dat_s1_translator_avalon_anti_slave_0_address;                                                 // sd_dat_s1_translator:av_address -> sd_dat:address
	wire          sd_dat_s1_translator_avalon_anti_slave_0_chipselect;                                              // sd_dat_s1_translator:av_chipselect -> sd_dat:chipselect
	wire          sd_dat_s1_translator_avalon_anti_slave_0_write;                                                   // sd_dat_s1_translator:av_write -> sd_dat:write_n
	wire   [31:0] sd_dat_s1_translator_avalon_anti_slave_0_readdata;                                                // sd_dat:readdata -> sd_dat_s1_translator:av_readdata
	wire    [1:0] sd_wp_n_s1_translator_avalon_anti_slave_0_address;                                                // sd_wp_n_s1_translator:av_address -> sd_wp_n:address
	wire   [31:0] sd_wp_n_s1_translator_avalon_anti_slave_0_readdata;                                               // sd_wp_n:readdata -> sd_wp_n_s1_translator:av_readdata
	wire   [31:0] epp_i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                          // epp_i2c_scl_s1_translator:av_writedata -> epp_i2c_scl:writedata
	wire    [1:0] epp_i2c_scl_s1_translator_avalon_anti_slave_0_address;                                            // epp_i2c_scl_s1_translator:av_address -> epp_i2c_scl:address
	wire          epp_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                         // epp_i2c_scl_s1_translator:av_chipselect -> epp_i2c_scl:chipselect
	wire          epp_i2c_scl_s1_translator_avalon_anti_slave_0_write;                                              // epp_i2c_scl_s1_translator:av_write -> epp_i2c_scl:write_n
	wire   [31:0] epp_i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                           // epp_i2c_scl:readdata -> epp_i2c_scl_s1_translator:av_readdata
	wire   [31:0] epp_i2c_sda_s1_translator_avalon_anti_slave_0_writedata;                                          // epp_i2c_sda_s1_translator:av_writedata -> epp_i2c_sda:writedata
	wire    [1:0] epp_i2c_sda_s1_translator_avalon_anti_slave_0_address;                                            // epp_i2c_sda_s1_translator:av_address -> epp_i2c_sda:address
	wire          epp_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect;                                         // epp_i2c_sda_s1_translator:av_chipselect -> epp_i2c_sda:chipselect
	wire          epp_i2c_sda_s1_translator_avalon_anti_slave_0_write;                                              // epp_i2c_sda_s1_translator:av_write -> epp_i2c_sda:write_n
	wire   [31:0] epp_i2c_sda_s1_translator_avalon_anti_slave_0_readdata;                                           // epp_i2c_sda:readdata -> epp_i2c_sda_s1_translator:av_readdata
	wire    [7:0] seg7_avalon_slave_translator_avalon_anti_slave_0_writedata;                                       // seg7_avalon_slave_translator:av_writedata -> seg7:s_writedata
	wire    [2:0] seg7_avalon_slave_translator_avalon_anti_slave_0_address;                                         // seg7_avalon_slave_translator:av_address -> seg7:s_address
	wire          seg7_avalon_slave_translator_avalon_anti_slave_0_write;                                           // seg7_avalon_slave_translator:av_write -> seg7:s_write
	wire          seg7_avalon_slave_translator_avalon_anti_slave_0_read;                                            // seg7_avalon_slave_translator:av_read -> seg7:s_read
	wire    [7:0] seg7_avalon_slave_translator_avalon_anti_slave_0_readdata;                                        // seg7:s_readdata -> seg7_avalon_slave_translator:av_readdata
	wire   [31:0] sw_s1_translator_avalon_anti_slave_0_writedata;                                                   // sw_s1_translator:av_writedata -> sw:writedata
	wire    [1:0] sw_s1_translator_avalon_anti_slave_0_address;                                                     // sw_s1_translator:av_address -> sw:address
	wire          sw_s1_translator_avalon_anti_slave_0_chipselect;                                                  // sw_s1_translator:av_chipselect -> sw:chipselect
	wire          sw_s1_translator_avalon_anti_slave_0_write;                                                       // sw_s1_translator:av_write -> sw:write_n
	wire   [31:0] sw_s1_translator_avalon_anti_slave_0_readdata;                                                    // sw:readdata -> sw_s1_translator:av_readdata
	wire   [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                              // i2c_scl_s1_translator:av_writedata -> i2c_scl:writedata
	wire    [1:0] i2c_scl_s1_translator_avalon_anti_slave_0_address;                                                // i2c_scl_s1_translator:av_address -> i2c_scl:address
	wire          i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                             // i2c_scl_s1_translator:av_chipselect -> i2c_scl:chipselect
	wire          i2c_scl_s1_translator_avalon_anti_slave_0_write;                                                  // i2c_scl_s1_translator:av_write -> i2c_scl:write_n
	wire   [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                               // i2c_scl:readdata -> i2c_scl_s1_translator:av_readdata
	wire   [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_writedata;                                              // i2c_sda_s1_translator:av_writedata -> i2c_sda:writedata
	wire    [1:0] i2c_sda_s1_translator_avalon_anti_slave_0_address;                                                // i2c_sda_s1_translator:av_address -> i2c_sda:address
	wire          i2c_sda_s1_translator_avalon_anti_slave_0_chipselect;                                             // i2c_sda_s1_translator:av_chipselect -> i2c_sda:chipselect
	wire          i2c_sda_s1_translator_avalon_anti_slave_0_write;                                                  // i2c_sda_s1_translator:av_write -> i2c_sda:write_n
	wire   [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_readdata;                                               // i2c_sda:readdata -> i2c_sda_s1_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                  // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                    // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer:readdata -> timer_s1_translator:av_readdata
	wire   [31:0] ledg_s1_translator_avalon_anti_slave_0_writedata;                                                 // ledg_s1_translator:av_writedata -> ledg:writedata
	wire    [1:0] ledg_s1_translator_avalon_anti_slave_0_address;                                                   // ledg_s1_translator:av_address -> ledg:address
	wire          ledg_s1_translator_avalon_anti_slave_0_chipselect;                                                // ledg_s1_translator:av_chipselect -> ledg:chipselect
	wire          ledg_s1_translator_avalon_anti_slave_0_write;                                                     // ledg_s1_translator:av_write -> ledg:write_n
	wire   [31:0] ledg_s1_translator_avalon_anti_slave_0_readdata;                                                  // ledg:readdata -> ledg_s1_translator:av_readdata
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_writedata;                                                 // ledr_s1_translator:av_writedata -> ledr:writedata
	wire    [1:0] ledr_s1_translator_avalon_anti_slave_0_address;                                                   // ledr_s1_translator:av_address -> ledr:address
	wire          ledr_s1_translator_avalon_anti_slave_0_chipselect;                                                // ledr_s1_translator:av_chipselect -> ledr:chipselect
	wire          ledr_s1_translator_avalon_anti_slave_0_write;                                                     // ledr_s1_translator:av_write -> ledr:write_n
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_readdata;                                                  // ledr:readdata -> ledr_s1_translator:av_readdata
	wire    [1:0] ir_s1_translator_avalon_anti_slave_0_address;                                                     // ir_s1_translator:av_address -> ir:address
	wire   [31:0] ir_s1_translator_avalon_anti_slave_0_readdata;                                                    // ir:readdata -> ir_s1_translator:av_readdata
	wire   [15:0] rs232_s1_translator_avalon_anti_slave_0_writedata;                                                // rs232_s1_translator:av_writedata -> rs232:writedata
	wire    [2:0] rs232_s1_translator_avalon_anti_slave_0_address;                                                  // rs232_s1_translator:av_address -> rs232:address
	wire          rs232_s1_translator_avalon_anti_slave_0_chipselect;                                               // rs232_s1_translator:av_chipselect -> rs232:chipselect
	wire          rs232_s1_translator_avalon_anti_slave_0_write;                                                    // rs232_s1_translator:av_write -> rs232:write_n
	wire          rs232_s1_translator_avalon_anti_slave_0_read;                                                     // rs232_s1_translator:av_read -> rs232:read_n
	wire   [15:0] rs232_s1_translator_avalon_anti_slave_0_readdata;                                                 // rs232:readdata -> rs232_s1_translator:av_readdata
	wire          rs232_s1_translator_avalon_anti_slave_0_begintransfer;                                            // rs232_s1_translator:av_begintransfer -> rs232:begintransfer
	wire          sysid_control_slave_translator_avalon_anti_slave_0_address;                                       // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                      // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                     // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                       // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                        // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                        // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount;                         // sgdma_tx_descriptor_read_translator:uav_burstcount -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata;                          // sgdma_tx_descriptor_read_translator:uav_writedata -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address;                            // sgdma_tx_descriptor_read_translator:uav_address -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock;                               // sgdma_tx_descriptor_read_translator:uav_lock -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write;                              // sgdma_tx_descriptor_read_translator:uav_write -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read;                               // sgdma_tx_descriptor_read_translator:uav_read -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata;                           // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_read_translator:uav_readdata
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                        // sgdma_tx_descriptor_read_translator:uav_debugaccess -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable;                         // sgdma_tx_descriptor_read_translator:uav_byteenable -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                      // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                       // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount;                        // sgdma_tx_descriptor_write_translator:uav_burstcount -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata;                         // sgdma_tx_descriptor_write_translator:uav_writedata -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address;                           // sgdma_tx_descriptor_write_translator:uav_address -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock;                              // sgdma_tx_descriptor_write_translator:uav_lock -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write;                             // sgdma_tx_descriptor_write_translator:uav_write -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read;                              // sgdma_tx_descriptor_write_translator:uav_read -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata;                          // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_write_translator:uav_readdata
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                       // sgdma_tx_descriptor_write_translator:uav_debugaccess -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable;                        // sgdma_tx_descriptor_write_translator:uav_byteenable -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                     // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                        // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount;                         // sgdma_rx_descriptor_read_translator:uav_burstcount -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata;                          // sgdma_rx_descriptor_read_translator:uav_writedata -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address;                            // sgdma_rx_descriptor_read_translator:uav_address -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock;                               // sgdma_rx_descriptor_read_translator:uav_lock -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write;                              // sgdma_rx_descriptor_read_translator:uav_write -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read;                               // sgdma_rx_descriptor_read_translator:uav_read -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata;                           // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_read_translator:uav_readdata
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                        // sgdma_rx_descriptor_read_translator:uav_debugaccess -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable;                         // sgdma_rx_descriptor_read_translator:uav_byteenable -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                      // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                       // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount;                        // sgdma_rx_descriptor_write_translator:uav_burstcount -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata;                         // sgdma_rx_descriptor_write_translator:uav_writedata -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address;                           // sgdma_rx_descriptor_write_translator:uav_address -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock;                              // sgdma_rx_descriptor_write_translator:uav_lock -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write;                             // sgdma_rx_descriptor_write_translator:uav_write -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read;                              // sgdma_rx_descriptor_write_translator:uav_read -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata;                          // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_write_translator:uav_readdata
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                       // sgdma_rx_descriptor_write_translator:uav_debugaccess -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable;                        // sgdma_rx_descriptor_write_translator:uav_byteenable -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                     // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest;                                 // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_m_read_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount;                                  // sgdma_tx_m_read_translator:uav_burstcount -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_writedata;                                   // sgdma_tx_m_read_translator:uav_writedata -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_address;                                     // sgdma_tx_m_read_translator:uav_address -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_lock;                                        // sgdma_tx_m_read_translator:uav_lock -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_write;                                       // sgdma_tx_m_read_translator:uav_write -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_read;                                        // sgdma_tx_m_read_translator:uav_read -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_readdata;                                    // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_m_read_translator:uav_readdata
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess;                                 // sgdma_tx_m_read_translator:uav_debugaccess -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable;                                  // sgdma_tx_m_read_translator:uav_byteenable -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid;                               // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_m_read_translator:uav_readdatavalid
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest;                                // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_m_write_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount;                                 // sgdma_rx_m_write_translator:uav_burstcount -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_writedata;                                  // sgdma_rx_m_write_translator:uav_writedata -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_address;                                    // sgdma_rx_m_write_translator:uav_address -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_lock;                                       // sgdma_rx_m_write_translator:uav_lock -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_write;                                      // sgdma_rx_m_write_translator:uav_write -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_read;                                       // sgdma_rx_m_write_translator:uav_read -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_readdata;                                   // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_m_write_translator:uav_readdata
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess;                                // sgdma_rx_m_write_translator:uav_debugaccess -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable;                                 // sgdma_rx_m_write_translator:uav_byteenable -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid;                              // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_m_write_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // cfi_flash_uas_translator:uav_waitrequest -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_uas_translator:uav_burstcount
	wire    [7:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                             // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_uas_translator:uav_writedata
	wire   [31:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_address;                               // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_uas_translator:uav_address
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_write;                                 // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_uas_translator:uav_write
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                  // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_uas_translator:uav_lock
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_read;                                  // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_uas_translator:uav_read
	wire    [7:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                              // cfi_flash_uas_translator:uav_readdata -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // cfi_flash_uas_translator:uav_readdatavalid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_uas_translator:uav_debugaccess
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_uas_translator:uav_byteenable
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                           // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // onchip_memory2_s1_translator:uav_waitrequest -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_s1_translator:uav_writedata
	wire   [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_s1_translator:uav_address
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_s1_translator:uav_write
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_s1_translator:uav_lock
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_s1_translator:uav_read
	wire   [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // onchip_memory2_s1_translator:uav_readdata -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // onchip_memory2_s1_translator:uav_readdatavalid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_s1_translator:uav_byteenable
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [3:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sram_avalon_slave_translator:uav_waitrequest -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_avalon_slave_translator:uav_burstcount
	wire   [15:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_avalon_slave_translator:uav_writedata
	wire   [31:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_avalon_slave_translator:uav_address
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_avalon_slave_translator:uav_write
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_avalon_slave_translator:uav_lock
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_avalon_slave_translator:uav_read
	wire   [15:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sram_avalon_slave_translator:uav_readdata -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sram_avalon_slave_translator:uav_readdatavalid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_avalon_slave_translator:uav_debugaccess
	wire    [1:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_avalon_slave_translator:uav_byteenable
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // clock_crossing_io_s0_translator:uav_waitrequest -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> clock_crossing_io_s0_translator:uav_burstcount
	wire   [31:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                      // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> clock_crossing_io_s0_translator:uav_writedata
	wire   [31:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_address;                        // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_address -> clock_crossing_io_s0_translator:uav_address
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_write;                          // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_write -> clock_crossing_io_s0_translator:uav_write
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_lock;                           // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_lock -> clock_crossing_io_s0_translator:uav_lock
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_read;                           // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_read -> clock_crossing_io_s0_translator:uav_read
	wire   [31:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                       // clock_crossing_io_s0_translator:uav_readdata -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // clock_crossing_io_s0_translator:uav_readdatavalid -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> clock_crossing_io_s0_translator:uav_debugaccess
	wire    [3:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> clock_crossing_io_s0_translator:uav_byteenable
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                    // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // audio_avalon_slave_translator:uav_waitrequest -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_avalon_slave_translator:uav_burstcount
	wire   [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_avalon_slave_translator:uav_writedata
	wire   [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_avalon_slave_translator:uav_address
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_avalon_slave_translator:uav_write
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_avalon_slave_translator:uav_lock
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_avalon_slave_translator:uav_read
	wire   [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // audio_avalon_slave_translator:uav_readdata -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // audio_avalon_slave_translator:uav_readdatavalid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_avalon_slave_translator:uav_debugaccess
	wire    [3:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_avalon_slave_translator:uav_byteenable
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // altpll_pll_slave_translator:uav_waitrequest -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_pll_slave_translator:uav_burstcount
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_pll_slave_translator:uav_writedata
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_pll_slave_translator:uav_address
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_pll_slave_translator:uav_write
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_pll_slave_translator:uav_lock
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_pll_slave_translator:uav_read
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // altpll_pll_slave_translator:uav_readdata -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // altpll_pll_slave_translator:uav_readdatavalid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_pll_slave_translator:uav_debugaccess
	wire    [3:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_pll_slave_translator:uav_byteenable
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // sma_in_s1_translator:uav_waitrequest -> sma_in_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sma_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sma_in_s1_translator:uav_burstcount
	wire   [31:0] sma_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sma_in_s1_translator:uav_writedata
	wire   [31:0] sma_in_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_address -> sma_in_s1_translator:uav_address
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_write -> sma_in_s1_translator:uav_write
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sma_in_s1_translator:uav_lock
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_read -> sma_in_s1_translator:uav_read
	wire   [31:0] sma_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // sma_in_s1_translator:uav_readdata -> sma_in_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // sma_in_s1_translator:uav_readdatavalid -> sma_in_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sma_in_s1_translator:uav_debugaccess
	wire    [3:0] sma_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // sma_in_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sma_in_s1_translator:uav_byteenable
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // sma_in_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // sma_in_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // sma_in_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // sma_in_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sma_in_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sma_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sma_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sma_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sma_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // sma_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // sma_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sma_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // sma_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sma_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // sma_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sma_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // sma_out_s1_translator:uav_waitrequest -> sma_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sma_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sma_out_s1_translator:uav_burstcount
	wire   [31:0] sma_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sma_out_s1_translator:uav_writedata
	wire   [31:0] sma_out_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> sma_out_s1_translator:uav_address
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> sma_out_s1_translator:uav_write
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sma_out_s1_translator:uav_lock
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> sma_out_s1_translator:uav_read
	wire   [31:0] sma_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // sma_out_s1_translator:uav_readdata -> sma_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // sma_out_s1_translator:uav_readdatavalid -> sma_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sma_out_s1_translator:uav_debugaccess
	wire    [3:0] sma_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // sma_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sma_out_s1_translator:uav_byteenable
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // sma_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // sma_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // sma_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // sma_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sma_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sma_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sma_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sma_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sma_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // sma_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // sma_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sma_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // sma_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sma_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // sma_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sma_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // ISP1362_IF_0_dc_translator:uav_waitrequest -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_burstcount -> ISP1362_IF_0_dc_translator:uav_burstcount
	wire   [31:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_writedata;                           // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_writedata -> ISP1362_IF_0_dc_translator:uav_writedata
	wire   [31:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_address;                             // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_address -> ISP1362_IF_0_dc_translator:uav_address
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_write;                               // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_write -> ISP1362_IF_0_dc_translator:uav_write
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_lock;                                // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_lock -> ISP1362_IF_0_dc_translator:uav_lock
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_read;                                // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_read -> ISP1362_IF_0_dc_translator:uav_read
	wire   [31:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_readdata;                            // ISP1362_IF_0_dc_translator:uav_readdata -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // ISP1362_IF_0_dc_translator:uav_readdatavalid -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ISP1362_IF_0_dc_translator:uav_debugaccess
	wire    [3:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:m0_byteenable -> ISP1362_IF_0_dc_translator:uav_byteenable
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_source_valid -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_data;                         // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_source_data -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // ISP1362_IF_0_hc_translator:uav_waitrequest -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_burstcount -> ISP1362_IF_0_hc_translator:uav_burstcount
	wire   [31:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_writedata;                           // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_writedata -> ISP1362_IF_0_hc_translator:uav_writedata
	wire   [31:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_address;                             // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_address -> ISP1362_IF_0_hc_translator:uav_address
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_write;                               // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_write -> ISP1362_IF_0_hc_translator:uav_write
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_lock;                                // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_lock -> ISP1362_IF_0_hc_translator:uav_lock
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_read;                                // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_read -> ISP1362_IF_0_hc_translator:uav_read
	wire   [31:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_readdata;                            // ISP1362_IF_0_hc_translator:uav_readdata -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // ISP1362_IF_0_hc_translator:uav_readdatavalid -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ISP1362_IF_0_hc_translator:uav_debugaccess
	wire    [3:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:m0_byteenable -> ISP1362_IF_0_hc_translator:uav_byteenable
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_source_valid -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_data;                         // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_source_data -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // descriptor_memory_s1_translator:uav_waitrequest -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_memory_s1_translator:uav_burstcount
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_memory_s1_translator:uav_writedata
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_memory_s1_translator:uav_address
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                          // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_memory_s1_translator:uav_write
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_memory_s1_translator:uav_lock
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_memory_s1_translator:uav_read
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                       // descriptor_memory_s1_translator:uav_readdata -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // descriptor_memory_s1_translator:uav_readdatavalid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_memory_s1_translator:uav_debugaccess
	wire    [3:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_memory_s1_translator:uav_byteenable
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // sgdma_rx_csr_translator:uav_waitrequest -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_rx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_rx_csr_translator:uav_writedata
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_rx_csr_translator:uav_address
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                  // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_rx_csr_translator:uav_write
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_rx_csr_translator:uav_lock
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_rx_csr_translator:uav_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                               // sgdma_rx_csr_translator:uav_readdata -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // sgdma_rx_csr_translator:uav_readdatavalid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_rx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_rx_csr_translator:uav_byteenable
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // sgdma_tx_csr_translator:uav_waitrequest -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_tx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_tx_csr_translator:uav_writedata
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_tx_csr_translator:uav_address
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                  // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_tx_csr_translator:uav_write
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_tx_csr_translator:uav_lock
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_tx_csr_translator:uav_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                               // sgdma_tx_csr_translator:uav_readdata -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // sgdma_tx_csr_translator:uav_readdatavalid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_tx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_tx_csr_translator:uav_byteenable
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // tse_mac_control_port_translator:uav_waitrequest -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_mac_control_port_translator:uav_burstcount
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_mac_control_port_translator:uav_writedata
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address;                        // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_address -> tse_mac_control_port_translator:uav_address
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write;                          // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_write -> tse_mac_control_port_translator:uav_write
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> tse_mac_control_port_translator:uav_lock
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read;                           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_read -> tse_mac_control_port_translator:uav_read
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                       // tse_mac_control_port_translator:uav_readdata -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // tse_mac_control_port_translator:uav_readdatavalid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_mac_control_port_translator:uav_debugaccess
	wire    [3:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_mac_control_port_translator:uav_byteenable
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // pio_0_s1_translator:uav_waitrequest -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_0_s1_translator:uav_burstcount
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_0_s1_translator:uav_writedata
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_0_s1_translator:uav_address
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_0_s1_translator:uav_write
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_0_s1_translator:uav_lock
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_0_s1_translator:uav_read
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // pio_0_s1_translator:uav_readdata -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // pio_0_s1_translator:uav_readdatavalid -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_0_s1_translator:uav_debugaccess
	wire    [3:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_0_s1_translator:uav_byteenable
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // pio_1_s1_translator:uav_waitrequest -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_1_s1_translator:uav_burstcount
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_1_s1_translator:uav_writedata
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_1_s1_translator:uav_address
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_1_s1_translator:uav_write
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_1_s1_translator:uav_lock
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_1_s1_translator:uav_read
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // pio_1_s1_translator:uav_readdata -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // pio_1_s1_translator:uav_readdatavalid -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_1_s1_translator:uav_debugaccess
	wire    [3:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_1_s1_translator:uav_byteenable
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_waitrequest;                            // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> clock_crossing_io_m0_translator:uav_waitrequest
	wire    [2:0] clock_crossing_io_m0_translator_avalon_universal_master_0_burstcount;                             // clock_crossing_io_m0_translator:uav_burstcount -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] clock_crossing_io_m0_translator_avalon_universal_master_0_writedata;                              // clock_crossing_io_m0_translator:uav_writedata -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [8:0] clock_crossing_io_m0_translator_avalon_universal_master_0_address;                                // clock_crossing_io_m0_translator:uav_address -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_address
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_lock;                                   // clock_crossing_io_m0_translator:uav_lock -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_write;                                  // clock_crossing_io_m0_translator:uav_write -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_write
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_read;                                   // clock_crossing_io_m0_translator:uav_read -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] clock_crossing_io_m0_translator_avalon_universal_master_0_readdata;                               // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_readdata -> clock_crossing_io_m0_translator:uav_readdata
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_debugaccess;                            // clock_crossing_io_m0_translator:uav_debugaccess -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] clock_crossing_io_m0_translator_avalon_universal_master_0_byteenable;                             // clock_crossing_io_m0_translator:uav_byteenable -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_readdatavalid;                          // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> clock_crossing_io_m0_translator:uav_readdatavalid
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // key_s1_translator:uav_waitrequest -> key_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // key_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key_s1_translator:uav_burstcount
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // key_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key_s1_translator:uav_writedata
	wire    [8:0] key_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // key_s1_translator_avalon_universal_slave_0_agent:m0_address -> key_s1_translator:uav_address
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // key_s1_translator_avalon_universal_slave_0_agent:m0_write -> key_s1_translator:uav_write
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // key_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key_s1_translator:uav_lock
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // key_s1_translator_avalon_universal_slave_0_agent:m0_read -> key_s1_translator:uav_read
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // key_s1_translator:uav_readdata -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // key_s1_translator:uav_readdatavalid -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // key_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key_s1_translator:uav_debugaccess
	wire    [3:0] key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // key_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key_s1_translator:uav_byteenable
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // key_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // key_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // key_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] key_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // key_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // key_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // lcd_control_slave_translator:uav_waitrequest -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_control_slave_translator:uav_burstcount
	wire   [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_control_slave_translator:uav_writedata
	wire    [8:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_control_slave_translator:uav_address
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_control_slave_translator:uav_write
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_control_slave_translator:uav_lock
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_control_slave_translator:uav_read
	wire   [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // lcd_control_slave_translator:uav_readdata -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // lcd_control_slave_translator:uav_readdatavalid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_control_slave_translator:uav_debugaccess
	wire    [3:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_control_slave_translator:uav_byteenable
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // sd_clk_s1_translator:uav_waitrequest -> sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_clk_s1_translator:uav_burstcount
	wire   [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_clk_s1_translator:uav_writedata
	wire    [8:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_address -> sd_clk_s1_translator:uav_address
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_write -> sd_clk_s1_translator:uav_write
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sd_clk_s1_translator:uav_lock
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_read -> sd_clk_s1_translator:uav_read
	wire   [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // sd_clk_s1_translator:uav_readdata -> sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // sd_clk_s1_translator:uav_readdatavalid -> sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_clk_s1_translator:uav_debugaccess
	wire    [3:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // sd_clk_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_clk_s1_translator:uav_byteenable
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // sd_clk_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // sd_clk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // sd_clk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // sd_clk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // sd_cmd_s1_translator:uav_waitrequest -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_cmd_s1_translator:uav_burstcount
	wire   [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_cmd_s1_translator:uav_writedata
	wire    [8:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_address -> sd_cmd_s1_translator:uav_address
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_write -> sd_cmd_s1_translator:uav_write
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sd_cmd_s1_translator:uav_lock
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_read -> sd_cmd_s1_translator:uav_read
	wire   [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // sd_cmd_s1_translator:uav_readdata -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // sd_cmd_s1_translator:uav_readdatavalid -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_cmd_s1_translator:uav_debugaccess
	wire    [3:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // sd_cmd_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_cmd_s1_translator:uav_byteenable
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // sd_dat_s1_translator:uav_waitrequest -> sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_dat_s1_translator:uav_burstcount
	wire   [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_dat_s1_translator:uav_writedata
	wire    [8:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_address -> sd_dat_s1_translator:uav_address
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_write -> sd_dat_s1_translator:uav_write
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sd_dat_s1_translator:uav_lock
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_read -> sd_dat_s1_translator:uav_read
	wire   [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // sd_dat_s1_translator:uav_readdata -> sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // sd_dat_s1_translator:uav_readdatavalid -> sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_dat_s1_translator:uav_debugaccess
	wire    [3:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // sd_dat_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_dat_s1_translator:uav_byteenable
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // sd_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // sd_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // sd_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // sd_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // sd_wp_n_s1_translator:uav_waitrequest -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_wp_n_s1_translator:uav_burstcount
	wire   [31:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_wp_n_s1_translator:uav_writedata
	wire    [8:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_address -> sd_wp_n_s1_translator:uav_address
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_write -> sd_wp_n_s1_translator:uav_write
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sd_wp_n_s1_translator:uav_lock
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_read -> sd_wp_n_s1_translator:uav_read
	wire   [31:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // sd_wp_n_s1_translator:uav_readdata -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // sd_wp_n_s1_translator:uav_readdatavalid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_wp_n_s1_translator:uav_debugaccess
	wire    [3:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_wp_n_s1_translator:uav_byteenable
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // epp_i2c_scl_s1_translator:uav_waitrequest -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> epp_i2c_scl_s1_translator:uav_burstcount
	wire   [31:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> epp_i2c_scl_s1_translator:uav_writedata
	wire    [8:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> epp_i2c_scl_s1_translator:uav_address
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> epp_i2c_scl_s1_translator:uav_write
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> epp_i2c_scl_s1_translator:uav_lock
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> epp_i2c_scl_s1_translator:uav_read
	wire   [31:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // epp_i2c_scl_s1_translator:uav_readdata -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // epp_i2c_scl_s1_translator:uav_readdatavalid -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epp_i2c_scl_s1_translator:uav_debugaccess
	wire    [3:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> epp_i2c_scl_s1_translator:uav_byteenable
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // epp_i2c_sda_s1_translator:uav_waitrequest -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> epp_i2c_sda_s1_translator:uav_burstcount
	wire   [31:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> epp_i2c_sda_s1_translator:uav_writedata
	wire    [8:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_address -> epp_i2c_sda_s1_translator:uav_address
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_write -> epp_i2c_sda_s1_translator:uav_write
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_lock -> epp_i2c_sda_s1_translator:uav_lock
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_read -> epp_i2c_sda_s1_translator:uav_read
	wire   [31:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // epp_i2c_sda_s1_translator:uav_readdata -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // epp_i2c_sda_s1_translator:uav_readdatavalid -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epp_i2c_sda_s1_translator:uav_debugaccess
	wire    [3:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> epp_i2c_sda_s1_translator:uav_byteenable
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // seg7_avalon_slave_translator:uav_waitrequest -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> seg7_avalon_slave_translator:uav_burstcount
	wire   [31:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> seg7_avalon_slave_translator:uav_writedata
	wire    [8:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> seg7_avalon_slave_translator:uav_address
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> seg7_avalon_slave_translator:uav_write
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> seg7_avalon_slave_translator:uav_lock
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> seg7_avalon_slave_translator:uav_read
	wire   [31:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // seg7_avalon_slave_translator:uav_readdata -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // seg7_avalon_slave_translator:uav_readdatavalid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seg7_avalon_slave_translator:uav_debugaccess
	wire    [3:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> seg7_avalon_slave_translator:uav_byteenable
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // sw_s1_translator:uav_waitrequest -> sw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // sw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sw_s1_translator:uav_burstcount
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // sw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sw_s1_translator:uav_writedata
	wire    [8:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // sw_s1_translator_avalon_universal_slave_0_agent:m0_address -> sw_s1_translator:uav_address
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // sw_s1_translator_avalon_universal_slave_0_agent:m0_write -> sw_s1_translator:uav_write
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // sw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sw_s1_translator:uav_lock
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // sw_s1_translator_avalon_universal_slave_0_agent:m0_read -> sw_s1_translator:uav_read
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // sw_s1_translator:uav_readdata -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // sw_s1_translator:uav_readdatavalid -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // sw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sw_s1_translator:uav_debugaccess
	wire    [3:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // sw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sw_s1_translator:uav_byteenable
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // i2c_scl_s1_translator:uav_waitrequest -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> i2c_scl_s1_translator:uav_burstcount
	wire   [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> i2c_scl_s1_translator:uav_writedata
	wire    [8:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> i2c_scl_s1_translator:uav_address
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> i2c_scl_s1_translator:uav_write
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> i2c_scl_s1_translator:uav_lock
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> i2c_scl_s1_translator:uav_read
	wire   [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // i2c_scl_s1_translator:uav_readdata -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // i2c_scl_s1_translator:uav_readdatavalid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> i2c_scl_s1_translator:uav_debugaccess
	wire    [3:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> i2c_scl_s1_translator:uav_byteenable
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // i2c_sda_s1_translator:uav_waitrequest -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> i2c_sda_s1_translator:uav_burstcount
	wire   [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> i2c_sda_s1_translator:uav_writedata
	wire    [8:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_address -> i2c_sda_s1_translator:uav_address
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_write -> i2c_sda_s1_translator:uav_write
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_lock -> i2c_sda_s1_translator:uav_lock
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_read -> i2c_sda_s1_translator:uav_read
	wire   [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // i2c_sda_s1_translator:uav_readdata -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // i2c_sda_s1_translator:uav_readdatavalid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> i2c_sda_s1_translator:uav_debugaccess
	wire    [3:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> i2c_sda_s1_translator:uav_byteenable
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire    [8:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // ledg_s1_translator:uav_waitrequest -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // ledg_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ledg_s1_translator:uav_burstcount
	wire   [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // ledg_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ledg_s1_translator:uav_writedata
	wire    [8:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // ledg_s1_translator_avalon_universal_slave_0_agent:m0_address -> ledg_s1_translator:uav_address
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // ledg_s1_translator_avalon_universal_slave_0_agent:m0_write -> ledg_s1_translator:uav_write
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // ledg_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ledg_s1_translator:uav_lock
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // ledg_s1_translator_avalon_universal_slave_0_agent:m0_read -> ledg_s1_translator:uav_read
	wire   [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // ledg_s1_translator:uav_readdata -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // ledg_s1_translator:uav_readdatavalid -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // ledg_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ledg_s1_translator:uav_debugaccess
	wire    [3:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // ledg_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ledg_s1_translator:uav_byteenable
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // ledr_s1_translator:uav_waitrequest -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // ledr_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ledr_s1_translator:uav_burstcount
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // ledr_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ledr_s1_translator:uav_writedata
	wire    [8:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // ledr_s1_translator_avalon_universal_slave_0_agent:m0_address -> ledr_s1_translator:uav_address
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // ledr_s1_translator_avalon_universal_slave_0_agent:m0_write -> ledr_s1_translator:uav_write
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // ledr_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ledr_s1_translator:uav_lock
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // ledr_s1_translator_avalon_universal_slave_0_agent:m0_read -> ledr_s1_translator:uav_read
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // ledr_s1_translator:uav_readdata -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // ledr_s1_translator:uav_readdatavalid -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // ledr_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ledr_s1_translator:uav_debugaccess
	wire    [3:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // ledr_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ledr_s1_translator:uav_byteenable
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // ir_s1_translator:uav_waitrequest -> ir_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // ir_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ir_s1_translator:uav_burstcount
	wire   [31:0] ir_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // ir_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ir_s1_translator:uav_writedata
	wire    [8:0] ir_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // ir_s1_translator_avalon_universal_slave_0_agent:m0_address -> ir_s1_translator:uav_address
	wire          ir_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // ir_s1_translator_avalon_universal_slave_0_agent:m0_write -> ir_s1_translator:uav_write
	wire          ir_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // ir_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ir_s1_translator:uav_lock
	wire          ir_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // ir_s1_translator_avalon_universal_slave_0_agent:m0_read -> ir_s1_translator:uav_read
	wire   [31:0] ir_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // ir_s1_translator:uav_readdata -> ir_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // ir_s1_translator:uav_readdatavalid -> ir_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // ir_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ir_s1_translator:uav_debugaccess
	wire    [3:0] ir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // ir_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ir_s1_translator:uav_byteenable
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // ir_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // ir_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // ir_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] ir_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // ir_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ir_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ir_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ir_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ir_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ir_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // ir_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // ir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // ir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // ir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // rs232_s1_translator:uav_waitrequest -> rs232_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // rs232_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> rs232_s1_translator:uav_burstcount
	wire   [31:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // rs232_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> rs232_s1_translator:uav_writedata
	wire    [8:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // rs232_s1_translator_avalon_universal_slave_0_agent:m0_address -> rs232_s1_translator:uav_address
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // rs232_s1_translator_avalon_universal_slave_0_agent:m0_write -> rs232_s1_translator:uav_write
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // rs232_s1_translator_avalon_universal_slave_0_agent:m0_lock -> rs232_s1_translator:uav_lock
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // rs232_s1_translator_avalon_universal_slave_0_agent:m0_read -> rs232_s1_translator:uav_read
	wire   [31:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // rs232_s1_translator:uav_readdata -> rs232_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // rs232_s1_translator:uav_readdatavalid -> rs232_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // rs232_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rs232_s1_translator:uav_debugaccess
	wire    [3:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // rs232_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> rs232_s1_translator:uav_byteenable
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // rs232_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // rs232_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // rs232_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // rs232_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rs232_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rs232_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rs232_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rs232_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rs232_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // rs232_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // rs232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rs232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // rs232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rs232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // rs232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rs232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire    [8:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [106:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [106:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;               // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                     // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;             // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [106:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                      // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_002:sink_ready -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;              // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                    // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;            // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [106:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                     // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                    // addr_router_003:sink_ready -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;               // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                     // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;             // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [106:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                      // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_004:sink_ready -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;              // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                    // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;            // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [106:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                     // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                    // addr_router_005:sink_ready -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid;                              // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire  [106:0] sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data;                               // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_006:sink_ready -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid;                             // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire  [106:0] sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data;                              // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_007:sink_ready -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [106:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                 // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [79:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_data;                                  // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_001:sink_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [106:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_002:sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [106:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_003:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [88:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_004:sink_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_valid;                          // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [106:0] clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_data;                           // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_005:sink_ready -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [106:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_007:sink_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [106:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_008:sink_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // sma_in_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // sma_in_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // sma_in_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [106:0] sma_in_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // sma_in_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          sma_in_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_009:sink_ready -> sma_in_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // sma_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // sma_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // sma_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [106:0] sma_out_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // sma_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          sma_out_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_010:sink_ready -> sma_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_valid;                               // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [106:0] isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_data;                                // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_011:sink_ready -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:rp_ready
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_valid;                               // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [106:0] isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_data;                                // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_012:sink_ready -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:rp_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                          // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [106:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_013:sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                  // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [106:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_014:sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                  // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [106:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_015:sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                          // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [106:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data;                           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_016:sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [106:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_017:sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [106:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_018:sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_valid;                         // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire   [83:0] clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_data;                          // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire          clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_008:sink_ready -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // key_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // key_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // key_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire   [83:0] key_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // key_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_019:sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire   [83:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_020:sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // sd_clk_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // sd_clk_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // sd_clk_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire   [83:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // sd_clk_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_021:sink_ready -> sd_clk_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire   [83:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // sd_cmd_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_022:sink_ready -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // sd_dat_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // sd_dat_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // sd_dat_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire   [83:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // sd_dat_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_023:sink_ready -> sd_dat_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire   [83:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_024:sink_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire   [83:0] epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_025:sink_ready -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire   [83:0] epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire          epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_026:sink_ready -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire   [83:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire          seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_027:sink_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // sw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // sw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // sw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire   [83:0] sw_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // sw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_028:sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire   [83:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_029:sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire   [83:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_030:sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire   [83:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_031:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // ledg_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // ledg_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // ledg_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire   [83:0] ledg_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // ledg_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_032:sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // ledr_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // ledr_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // ledr_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire   [83:0] ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // ledr_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_033:sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // ir_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // ir_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // ir_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire   [83:0] ir_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // ir_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire          ir_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_034:sink_ready -> ir_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // rs232_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // rs232_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // rs232_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire   [83:0] rs232_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // rs232_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire          rs232_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_035:sink_ready -> rs232_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire   [83:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_036:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                            // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [106:0] addr_router_src_data;                                                                             // addr_router:src_data -> limiter:cmd_sink_data
	wire   [18:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                            // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                      // limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                            // limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                    // limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_rsp_src_data;                                                                             // limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_rsp_src_channel;                                                                          // limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                            // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [106:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [18:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                        // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                  // limiter_001:rsp_src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                        // limiter_001:rsp_src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                // limiter_001:rsp_src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_001_rsp_src_data;                                                                         // limiter_001:rsp_src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_001_rsp_src_channel;                                                                      // limiter_001:rsp_src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                        // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_008_src_endofpacket;                                                                  // addr_router_008:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_008_src_valid;                                                                        // addr_router_008:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_008_src_startofpacket;                                                                // addr_router_008:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire   [83:0] addr_router_008_src_data;                                                                         // addr_router_008:src_data -> limiter_002:cmd_sink_data
	wire   [17:0] addr_router_008_src_channel;                                                                      // addr_router_008:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_008_src_ready;                                                                        // limiter_002:cmd_sink_ready -> addr_router_008:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                  // limiter_002:rsp_src_endofpacket -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                        // limiter_002:rsp_src_valid -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                // limiter_002:rsp_src_startofpacket -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [83:0] limiter_002_rsp_src_data;                                                                         // limiter_002:rsp_src_data -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [17:0] limiter_002_rsp_src_channel;                                                                      // limiter_002:rsp_src_channel -> clock_crossing_io_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                        // clock_crossing_io_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                // burst_adapter:source0_endofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                      // burst_adapter:source0_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                              // burst_adapter:source0_startofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_source0_data;                                                                       // burst_adapter:source0_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                      // cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [18:0] burst_adapter_source0_channel;                                                                    // burst_adapter:source0_channel -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                            // burst_adapter_001:source0_endofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                  // burst_adapter_001:source0_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                          // burst_adapter_001:source0_startofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_001_source0_data;                                                                   // burst_adapter_001:source0_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                  // sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [18:0] burst_adapter_001_source0_channel;                                                                // burst_adapter_001:source0_channel -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> [addr_router_008:reset, clock_crossing_io:m0_reset, clock_crossing_io_m0_translator:reset, clock_crossing_io_m0_translator_avalon_universal_master_0_agent:reset, cmd_xbar_demux_008:reset, epp_i2c_sda:reset_n, epp_i2c_sda_s1_translator:reset, epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:reset, epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, i2c_scl:reset_n, i2c_scl_s1_translator:reset, i2c_scl_s1_translator_avalon_universal_slave_0_agent:reset, i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, i2c_sda:reset_n, i2c_sda_s1_translator:reset, i2c_sda_s1_translator_avalon_universal_slave_0_agent:reset, i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, id_router_030:reset, id_router_031:reset, id_router_032:reset, id_router_033:reset, id_router_035:reset, id_router_036:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, key:reset_n, key_s1_translator:reset, key_s1_translator_avalon_universal_slave_0_agent:reset, key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd:reset_n, lcd_control_slave_translator:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ledg:reset_n, ledg_s1_translator:reset, ledg_s1_translator_avalon_universal_slave_0_agent:reset, ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ledr:reset_n, ledr_s1_translator:reset, ledr_s1_translator_avalon_universal_slave_0_agent:reset, ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_002:reset, rs232:reset_n, rs232_s1_translator:reset, rs232_s1_translator_avalon_universal_slave_0_agent:reset, rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_032:reset, rsp_xbar_demux_033:reset, rsp_xbar_demux_035:reset, rsp_xbar_demux_036:reset, rsp_xbar_mux_008:reset, sd_clk:reset_n, sd_clk_s1_translator:reset, sd_clk_s1_translator_avalon_universal_slave_0_agent:reset, sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sd_cmd:reset_n, sd_cmd_s1_translator:reset, sd_cmd_s1_translator_avalon_universal_slave_0_agent:reset, sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sd_dat:reset_n, sd_dat_s1_translator:reset, sd_dat_s1_translator_avalon_universal_slave_0_agent:reset, sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sd_wp_n:reset_n, sd_wp_n_s1_translator:reset, sd_wp_n_s1_translator_avalon_universal_slave_0_agent:reset, sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, seg7:s_reset, seg7_avalon_slave_translator:reset, seg7_avalon_slave_translator_avalon_universal_slave_0_agent:reset, seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sw:reset_n, sw_s1_translator:reset, sw_s1_translator_avalon_universal_slave_0_agent:reset, sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_001_reset_out_reset;                                                               // rst_controller_001:reset_out -> [ISP1362_IF_0:avs_hc_reset_n_iRST_N, ISP1362_IF_0_hc_translator:reset, ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:reset, ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, addr_router_006:reset, addr_router_007:reset, audio:avs_s1_reset, audio_avalon_slave_translator:reset, audio_avalon_slave_translator_avalon_universal_slave_0_agent:reset, audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter:reset, burst_adapter_001:reset, cfi_flash:reset_reset, cfi_flash_uas_translator:reset, cfi_flash_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, clock_crossing_io:s0_reset, clock_crossing_io_s0_translator:reset, clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:reset, clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_013:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, descriptor_memory:reset, descriptor_memory_s1_translator:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_009:reset, id_router_010:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, onchip_memory2:reset, onchip_memory2_s1_translator:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx:system_reset_n, sgdma_rx_csr_translator:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx_descriptor_read_translator:reset, sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_rx_descriptor_write_translator:reset, sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_rx_m_write_translator:reset, sgdma_rx_m_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx:system_reset_n, sgdma_tx_csr_translator:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_tx_descriptor_read_translator:reset, sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_tx_descriptor_write_translator:reset, sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx_m_read_translator:reset, sgdma_tx_m_read_translator_avalon_universal_master_0_agent:reset, sma_in:reset_n, sma_in_s1_translator:reset, sma_in_s1_translator_avalon_universal_slave_0_agent:reset, sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sma_out:reset_n, sma_out_s1_translator:reset, sma_out_s1_translator_avalon_universal_slave_0_agent:reset, sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram:reset_n, sram_avalon_slave_translator:reset, sram_avalon_slave_translator_avalon_universal_slave_0_agent:reset, sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tri_state_bridge_flash_bridge_0:reset, tri_state_flash_bridge_pinSharer_0:reset_reset, tse_mac:reset, tse_mac_control_port_translator:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_002_reset_out_reset;                                                               // rst_controller_002:reset_out -> [epp_i2c_scl:reset_n, epp_i2c_scl_s1_translator:reset, epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:reset, epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_025:reset, rsp_xbar_demux_025:reset]
	wire          rst_controller_003_reset_out_reset;                                                               // rst_controller_003:reset_out -> [altpll:reset, altpll_pll_slave_translator:reset, altpll_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_003:in_reset, id_router_008:reset, rsp_xbar_demux_008:reset]
	wire          rst_controller_004_reset_out_reset;                                                               // rst_controller_004:reset_out -> [id_router_034:reset, ir:reset_n, ir_s1_translator:reset, ir_s1_translator_avalon_universal_slave_0_agent:reset, ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_034:reset]
	wire          rst_controller_005_reset_out_reset;                                                               // rst_controller_005:reset_out -> [crosser_001:out_reset, crosser_002:out_reset, crosser_004:in_reset, crosser_005:in_reset, id_router_017:reset, id_router_018:reset, pio_0:reset_n, pio_0_s1_translator:reset, pio_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_1:reset_n, pio_1_s1_translator:reset, pio_1_s1_translator_avalon_universal_slave_0_agent:reset, pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [18:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [18:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [18:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                        // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                  // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                        // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src3_data;                                                                         // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [18:0] cmd_xbar_demux_src3_channel;                                                                      // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                        // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_src4_endofpacket;                                                                  // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                        // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src4_data;                                                                         // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [18:0] cmd_xbar_demux_src4_channel;                                                                      // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_src4_ready;                                                                        // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src1_data;                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src1_channel;                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                              // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                    // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                            // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src2_data;                                                                     // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src2_channel;                                                                  // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                    // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                              // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                    // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                            // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src3_data;                                                                     // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src3_channel;                                                                  // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                    // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                              // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                    // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                            // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src4_data;                                                                     // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src4_channel;                                                                  // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                    // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                              // cmd_xbar_demux_001:src5_endofpacket -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                    // cmd_xbar_demux_001:src5_valid -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                            // cmd_xbar_demux_001:src5_startofpacket -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src5_data;                                                                     // cmd_xbar_demux_001:src5_data -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src5_channel;                                                                  // cmd_xbar_demux_001:src5_channel -> clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                              // cmd_xbar_demux_001:src6_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                    // cmd_xbar_demux_001:src6_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                            // cmd_xbar_demux_001:src6_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src6_data;                                                                     // cmd_xbar_demux_001:src6_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src6_channel;                                                                  // cmd_xbar_demux_001:src6_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                              // cmd_xbar_demux_001:src7_endofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                    // cmd_xbar_demux_001:src7_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                            // cmd_xbar_demux_001:src7_startofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src7_data;                                                                     // cmd_xbar_demux_001:src7_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src7_channel;                                                                  // cmd_xbar_demux_001:src7_channel -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                              // cmd_xbar_demux_001:src9_endofpacket -> sma_in_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                    // cmd_xbar_demux_001:src9_valid -> sma_in_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                            // cmd_xbar_demux_001:src9_startofpacket -> sma_in_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src9_data;                                                                     // cmd_xbar_demux_001:src9_data -> sma_in_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src9_channel;                                                                  // cmd_xbar_demux_001:src9_channel -> sma_in_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                             // cmd_xbar_demux_001:src10_endofpacket -> sma_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                   // cmd_xbar_demux_001:src10_valid -> sma_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                           // cmd_xbar_demux_001:src10_startofpacket -> sma_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src10_data;                                                                    // cmd_xbar_demux_001:src10_data -> sma_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src10_channel;                                                                 // cmd_xbar_demux_001:src10_channel -> sma_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                             // cmd_xbar_demux_001:src11_endofpacket -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                   // cmd_xbar_demux_001:src11_valid -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                           // cmd_xbar_demux_001:src11_startofpacket -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src11_data;                                                                    // cmd_xbar_demux_001:src11_data -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src11_channel;                                                                 // cmd_xbar_demux_001:src11_channel -> ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                             // cmd_xbar_demux_001:src12_endofpacket -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                   // cmd_xbar_demux_001:src12_valid -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                           // cmd_xbar_demux_001:src12_startofpacket -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src12_data;                                                                    // cmd_xbar_demux_001:src12_data -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src12_channel;                                                                 // cmd_xbar_demux_001:src12_channel -> ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                             // cmd_xbar_demux_001:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                   // cmd_xbar_demux_001:src13_valid -> cmd_xbar_mux_013:sink0_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                           // cmd_xbar_demux_001:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src13_data;                                                                    // cmd_xbar_demux_001:src13_data -> cmd_xbar_mux_013:sink0_data
	wire   [18:0] cmd_xbar_demux_001_src13_channel;                                                                 // cmd_xbar_demux_001:src13_channel -> cmd_xbar_mux_013:sink0_channel
	wire          cmd_xbar_demux_001_src13_ready;                                                                   // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux_001:src13_ready
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                             // cmd_xbar_demux_001:src14_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                   // cmd_xbar_demux_001:src14_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                           // cmd_xbar_demux_001:src14_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src14_data;                                                                    // cmd_xbar_demux_001:src14_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src14_channel;                                                                 // cmd_xbar_demux_001:src14_channel -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                             // cmd_xbar_demux_001:src15_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                   // cmd_xbar_demux_001:src15_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                           // cmd_xbar_demux_001:src15_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src15_data;                                                                    // cmd_xbar_demux_001:src15_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src15_channel;                                                                 // cmd_xbar_demux_001:src15_channel -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                             // cmd_xbar_demux_001:src16_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                   // cmd_xbar_demux_001:src16_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                           // cmd_xbar_demux_001:src16_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src16_data;                                                                    // cmd_xbar_demux_001:src16_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src16_channel;                                                                 // cmd_xbar_demux_001:src16_channel -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                              // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                    // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_013:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                            // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src0_data;                                                                     // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_013:sink1_data
	wire   [18:0] cmd_xbar_demux_002_src0_channel;                                                                  // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_013:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                    // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                              // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_013:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                    // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_013:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                            // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_013:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src0_data;                                                                     // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_013:sink2_data
	wire   [18:0] cmd_xbar_demux_003_src0_channel;                                                                  // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_013:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                    // cmd_xbar_mux_013:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                              // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_013:sink3_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                    // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_013:sink3_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                            // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_013:sink3_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src0_data;                                                                     // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_013:sink3_data
	wire   [18:0] cmd_xbar_demux_004_src0_channel;                                                                  // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_013:sink3_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                    // cmd_xbar_mux_013:sink3_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                              // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_013:sink4_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                    // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_013:sink4_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                            // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_013:sink4_startofpacket
	wire  [106:0] cmd_xbar_demux_005_src0_data;                                                                     // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_013:sink4_data
	wire   [18:0] cmd_xbar_demux_005_src0_channel;                                                                  // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_013:sink4_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                    // cmd_xbar_mux_013:sink4_ready -> cmd_xbar_demux_005:src0_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                              // cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                    // cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_003:sink2_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                            // cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src0_data;                                                                     // cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_003:sink2_data
	wire   [18:0] cmd_xbar_demux_006_src0_channel;                                                                  // cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_003:sink2_channel
	wire          cmd_xbar_demux_006_src0_ready;                                                                    // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_006:src0_ready
	wire          cmd_xbar_demux_007_src0_endofpacket;                                                              // cmd_xbar_demux_007:src0_endofpacket -> cmd_xbar_mux_003:sink3_endofpacket
	wire          cmd_xbar_demux_007_src0_valid;                                                                    // cmd_xbar_demux_007:src0_valid -> cmd_xbar_mux_003:sink3_valid
	wire          cmd_xbar_demux_007_src0_startofpacket;                                                            // cmd_xbar_demux_007:src0_startofpacket -> cmd_xbar_mux_003:sink3_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src0_data;                                                                     // cmd_xbar_demux_007:src0_data -> cmd_xbar_mux_003:sink3_data
	wire   [18:0] cmd_xbar_demux_007_src0_channel;                                                                  // cmd_xbar_demux_007:src0_channel -> cmd_xbar_mux_003:sink3_channel
	wire          cmd_xbar_demux_007_src0_ready;                                                                    // cmd_xbar_mux_003:sink3_ready -> cmd_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [18:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [18:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                        // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [18:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src1_data;                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [18:0] rsp_xbar_demux_001_src1_channel;                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [18:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                              // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                    // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                            // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src1_data;                                                                     // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [18:0] rsp_xbar_demux_002_src1_channel;                                                                  // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                    // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [18:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                    // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                              // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                    // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                            // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src1_data;                                                                     // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [18:0] rsp_xbar_demux_003_src1_channel;                                                                  // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                    // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_003_src2_endofpacket;                                                              // rsp_xbar_demux_003:src2_endofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src2_valid;                                                                    // rsp_xbar_demux_003:src2_valid -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src2_startofpacket;                                                            // rsp_xbar_demux_003:src2_startofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src2_data;                                                                     // rsp_xbar_demux_003:src2_data -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] rsp_xbar_demux_003_src2_channel;                                                                  // rsp_xbar_demux_003:src2_channel -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src3_endofpacket;                                                              // rsp_xbar_demux_003:src3_endofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src3_valid;                                                                    // rsp_xbar_demux_003:src3_valid -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src3_startofpacket;                                                            // rsp_xbar_demux_003:src3_startofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src3_data;                                                                     // rsp_xbar_demux_003:src3_data -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] rsp_xbar_demux_003_src3_channel;                                                                  // rsp_xbar_demux_003:src3_channel -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                              // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                    // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                            // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                     // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [18:0] rsp_xbar_demux_004_src0_channel;                                                                  // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                    // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                              // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                    // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                            // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src1_data;                                                                     // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [18:0] rsp_xbar_demux_004_src1_channel;                                                                  // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                    // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                              // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                    // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                            // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src0_data;                                                                     // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [18:0] rsp_xbar_demux_005_src0_channel;                                                                  // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                    // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                              // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                    // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                            // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                     // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [18:0] rsp_xbar_demux_006_src0_channel;                                                                  // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                    // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                              // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                    // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                            // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_007_src0_data;                                                                     // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [18:0] rsp_xbar_demux_007_src0_channel;                                                                  // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                    // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                              // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                    // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                            // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src0_data;                                                                     // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [18:0] rsp_xbar_demux_009_src0_channel;                                                                  // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                    // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                              // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                    // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                            // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src0_data;                                                                     // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [18:0] rsp_xbar_demux_010_src0_channel;                                                                  // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                    // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                              // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                    // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                            // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [106:0] rsp_xbar_demux_011_src0_data;                                                                     // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [18:0] rsp_xbar_demux_011_src0_channel;                                                                  // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                    // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                              // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                    // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                            // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [106:0] rsp_xbar_demux_012_src0_data;                                                                     // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [18:0] rsp_xbar_demux_012_src0_channel;                                                                  // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                    // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                              // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                    // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                            // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src0_data;                                                                     // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [18:0] rsp_xbar_demux_013_src0_channel;                                                                  // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                    // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_013_src1_endofpacket;                                                              // rsp_xbar_demux_013:src1_endofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_013_src1_valid;                                                                    // rsp_xbar_demux_013:src1_valid -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_013_src1_startofpacket;                                                            // rsp_xbar_demux_013:src1_startofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src1_data;                                                                     // rsp_xbar_demux_013:src1_data -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] rsp_xbar_demux_013_src1_channel;                                                                  // rsp_xbar_demux_013:src1_channel -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_013_src2_endofpacket;                                                              // rsp_xbar_demux_013:src2_endofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_013_src2_valid;                                                                    // rsp_xbar_demux_013:src2_valid -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_013_src2_startofpacket;                                                            // rsp_xbar_demux_013:src2_startofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src2_data;                                                                     // rsp_xbar_demux_013:src2_data -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] rsp_xbar_demux_013_src2_channel;                                                                  // rsp_xbar_demux_013:src2_channel -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_013_src3_endofpacket;                                                              // rsp_xbar_demux_013:src3_endofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_013_src3_valid;                                                                    // rsp_xbar_demux_013:src3_valid -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_013_src3_startofpacket;                                                            // rsp_xbar_demux_013:src3_startofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src3_data;                                                                     // rsp_xbar_demux_013:src3_data -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] rsp_xbar_demux_013_src3_channel;                                                                  // rsp_xbar_demux_013:src3_channel -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_013_src4_endofpacket;                                                              // rsp_xbar_demux_013:src4_endofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_013_src4_valid;                                                                    // rsp_xbar_demux_013:src4_valid -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_013_src4_startofpacket;                                                            // rsp_xbar_demux_013:src4_startofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src4_data;                                                                     // rsp_xbar_demux_013:src4_data -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] rsp_xbar_demux_013_src4_channel;                                                                  // rsp_xbar_demux_013:src4_channel -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                              // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                    // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                            // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [106:0] rsp_xbar_demux_014_src0_data;                                                                     // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [18:0] rsp_xbar_demux_014_src0_channel;                                                                  // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                    // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                              // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                    // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                            // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src0_data;                                                                     // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [18:0] rsp_xbar_demux_015_src0_channel;                                                                  // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                    // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                              // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                    // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                            // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [106:0] rsp_xbar_demux_016_src0_data;                                                                     // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [18:0] rsp_xbar_demux_016_src0_channel;                                                                  // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                    // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                      // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                    // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [106:0] limiter_cmd_src_data;                                                                             // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [18:0] limiter_cmd_src_channel;                                                                          // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                           // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                  // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [106:0] limiter_001_cmd_src_data;                                                                         // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [18:0] limiter_001_cmd_src_channel;                                                                      // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                 // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                       // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                               // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_001_src_data;                                                                        // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_001_src_channel;                                                                     // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                       // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                  // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                        // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [106:0] addr_router_002_src_data;                                                                         // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [18:0] addr_router_002_src_channel;                                                                      // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                        // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_013_src1_ready;                                                                    // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src1_ready
	wire          addr_router_003_src_endofpacket;                                                                  // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                        // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [106:0] addr_router_003_src_data;                                                                         // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [18:0] addr_router_003_src_channel;                                                                      // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                        // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_013_src2_ready;                                                                    // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src2_ready
	wire          addr_router_004_src_endofpacket;                                                                  // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                        // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [106:0] addr_router_004_src_data;                                                                         // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [18:0] addr_router_004_src_channel;                                                                      // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                        // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_013_src3_ready;                                                                    // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src3_ready
	wire          addr_router_005_src_endofpacket;                                                                  // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                        // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [106:0] addr_router_005_src_data;                                                                         // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire   [18:0] addr_router_005_src_channel;                                                                      // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                        // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          rsp_xbar_demux_013_src4_ready;                                                                    // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src4_ready
	wire          addr_router_006_src_endofpacket;                                                                  // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          addr_router_006_src_valid;                                                                        // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire          addr_router_006_src_startofpacket;                                                                // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire  [106:0] addr_router_006_src_data;                                                                         // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire   [18:0] addr_router_006_src_channel;                                                                      // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire          addr_router_006_src_ready;                                                                        // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire          rsp_xbar_demux_003_src2_ready;                                                                    // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src2_ready
	wire          addr_router_007_src_endofpacket;                                                                  // addr_router_007:src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire          addr_router_007_src_valid;                                                                        // addr_router_007:src_valid -> cmd_xbar_demux_007:sink_valid
	wire          addr_router_007_src_startofpacket;                                                                // addr_router_007:src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire  [106:0] addr_router_007_src_data;                                                                         // addr_router_007:src_data -> cmd_xbar_demux_007:sink_data
	wire   [18:0] addr_router_007_src_channel;                                                                      // addr_router_007:src_channel -> cmd_xbar_demux_007:sink_channel
	wire          addr_router_007_src_ready;                                                                        // cmd_xbar_demux_007:sink_ready -> addr_router_007:src_ready
	wire          rsp_xbar_demux_003_src3_ready;                                                                    // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src3_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [106:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [18:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                 // cmd_xbar_mux_002:src_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                       // cmd_xbar_mux_002:src_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                               // cmd_xbar_mux_002:src_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_002_src_data;                                                                        // cmd_xbar_mux_002:src_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_002_src_channel;                                                                     // cmd_xbar_mux_002:src_channel -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                          // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [106:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [18:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                          // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                 // cmd_xbar_mux_003:src_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                       // cmd_xbar_mux_003:src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                               // cmd_xbar_mux_003:src_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_003_src_data;                                                                        // cmd_xbar_mux_003:src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_003_src_channel;                                                                     // cmd_xbar_mux_003:src_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                       // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [106:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [18:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                    // clock_crossing_io_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [106:0] id_router_005_src_data;                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [18:0] id_router_005_src_channel;                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [18:0] id_router_006_src_channel;                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                    // audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                    // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                          // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                  // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [106:0] id_router_007_src_data;                                                                           // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [18:0] id_router_007_src_channel;                                                                        // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                          // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          crosser_out_ready;                                                                                // altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_008_src_endofpacket;                                                                    // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                          // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                  // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [106:0] id_router_008_src_data;                                                                           // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [18:0] id_router_008_src_channel;                                                                        // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                          // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                    // sma_in_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                    // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                          // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                  // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [106:0] id_router_009_src_data;                                                                           // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [18:0] id_router_009_src_channel;                                                                        // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                          // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                   // sma_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                    // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                          // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                  // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [106:0] id_router_010_src_data;                                                                           // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [18:0] id_router_010_src_channel;                                                                        // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                          // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                   // ISP1362_IF_0_dc_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                    // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                          // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                  // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [106:0] id_router_011_src_data;                                                                           // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [18:0] id_router_011_src_channel;                                                                        // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                          // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                   // ISP1362_IF_0_hc_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                    // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                          // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                  // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [106:0] id_router_012_src_data;                                                                           // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [18:0] id_router_012_src_channel;                                                                        // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                          // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_mux_013_src_endofpacket;                                                                 // cmd_xbar_mux_013:src_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_013_src_valid;                                                                       // cmd_xbar_mux_013:src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_013_src_startofpacket;                                                               // cmd_xbar_mux_013:src_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_013_src_data;                                                                        // cmd_xbar_mux_013:src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_013_src_channel;                                                                     // cmd_xbar_mux_013:src_channel -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_013_src_ready;                                                                       // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire          id_router_013_src_endofpacket;                                                                    // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                          // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                  // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [106:0] id_router_013_src_data;                                                                           // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [18:0] id_router_013_src_channel;                                                                        // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                          // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                    // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                          // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                  // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [106:0] id_router_014_src_data;                                                                           // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [18:0] id_router_014_src_channel;                                                                        // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                          // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                    // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                          // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                  // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [106:0] id_router_015_src_data;                                                                           // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [18:0] id_router_015_src_channel;                                                                        // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                          // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_001_src16_ready;                                                                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire          id_router_016_src_endofpacket;                                                                    // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                          // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                  // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [106:0] id_router_016_src_data;                                                                           // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [18:0] id_router_016_src_channel;                                                                        // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                          // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          crosser_001_out_ready;                                                                            // pio_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire          id_router_017_src_endofpacket;                                                                    // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                          // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                  // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [106:0] id_router_017_src_data;                                                                           // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [18:0] id_router_017_src_channel;                                                                        // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                          // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          crosser_002_out_ready;                                                                            // pio_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire          id_router_018_src_endofpacket;                                                                    // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                          // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                  // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [106:0] id_router_018_src_data;                                                                           // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [18:0] id_router_018_src_channel;                                                                        // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                          // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_008_src0_endofpacket;                                                              // cmd_xbar_demux_008:src0_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src0_valid;                                                                    // cmd_xbar_demux_008:src0_valid -> key_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src0_startofpacket;                                                            // cmd_xbar_demux_008:src0_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src0_data;                                                                     // cmd_xbar_demux_008:src0_data -> key_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src0_channel;                                                                  // cmd_xbar_demux_008:src0_channel -> key_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src1_endofpacket;                                                              // cmd_xbar_demux_008:src1_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src1_valid;                                                                    // cmd_xbar_demux_008:src1_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src1_startofpacket;                                                            // cmd_xbar_demux_008:src1_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src1_data;                                                                     // cmd_xbar_demux_008:src1_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src1_channel;                                                                  // cmd_xbar_demux_008:src1_channel -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src2_endofpacket;                                                              // cmd_xbar_demux_008:src2_endofpacket -> sd_clk_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src2_valid;                                                                    // cmd_xbar_demux_008:src2_valid -> sd_clk_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src2_startofpacket;                                                            // cmd_xbar_demux_008:src2_startofpacket -> sd_clk_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src2_data;                                                                     // cmd_xbar_demux_008:src2_data -> sd_clk_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src2_channel;                                                                  // cmd_xbar_demux_008:src2_channel -> sd_clk_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src3_endofpacket;                                                              // cmd_xbar_demux_008:src3_endofpacket -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src3_valid;                                                                    // cmd_xbar_demux_008:src3_valid -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src3_startofpacket;                                                            // cmd_xbar_demux_008:src3_startofpacket -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src3_data;                                                                     // cmd_xbar_demux_008:src3_data -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src3_channel;                                                                  // cmd_xbar_demux_008:src3_channel -> sd_cmd_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src4_endofpacket;                                                              // cmd_xbar_demux_008:src4_endofpacket -> sd_dat_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src4_valid;                                                                    // cmd_xbar_demux_008:src4_valid -> sd_dat_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src4_startofpacket;                                                            // cmd_xbar_demux_008:src4_startofpacket -> sd_dat_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src4_data;                                                                     // cmd_xbar_demux_008:src4_data -> sd_dat_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src4_channel;                                                                  // cmd_xbar_demux_008:src4_channel -> sd_dat_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src5_endofpacket;                                                              // cmd_xbar_demux_008:src5_endofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src5_valid;                                                                    // cmd_xbar_demux_008:src5_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src5_startofpacket;                                                            // cmd_xbar_demux_008:src5_startofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src5_data;                                                                     // cmd_xbar_demux_008:src5_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src5_channel;                                                                  // cmd_xbar_demux_008:src5_channel -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src6_endofpacket;                                                              // cmd_xbar_demux_008:src6_endofpacket -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src6_valid;                                                                    // cmd_xbar_demux_008:src6_valid -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src6_startofpacket;                                                            // cmd_xbar_demux_008:src6_startofpacket -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src6_data;                                                                     // cmd_xbar_demux_008:src6_data -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src6_channel;                                                                  // cmd_xbar_demux_008:src6_channel -> epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src7_endofpacket;                                                              // cmd_xbar_demux_008:src7_endofpacket -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src7_valid;                                                                    // cmd_xbar_demux_008:src7_valid -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src7_startofpacket;                                                            // cmd_xbar_demux_008:src7_startofpacket -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src7_data;                                                                     // cmd_xbar_demux_008:src7_data -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src7_channel;                                                                  // cmd_xbar_demux_008:src7_channel -> epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src8_endofpacket;                                                              // cmd_xbar_demux_008:src8_endofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src8_valid;                                                                    // cmd_xbar_demux_008:src8_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src8_startofpacket;                                                            // cmd_xbar_demux_008:src8_startofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src8_data;                                                                     // cmd_xbar_demux_008:src8_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src8_channel;                                                                  // cmd_xbar_demux_008:src8_channel -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src9_endofpacket;                                                              // cmd_xbar_demux_008:src9_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src9_valid;                                                                    // cmd_xbar_demux_008:src9_valid -> sw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src9_startofpacket;                                                            // cmd_xbar_demux_008:src9_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src9_data;                                                                     // cmd_xbar_demux_008:src9_data -> sw_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src9_channel;                                                                  // cmd_xbar_demux_008:src9_channel -> sw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src10_endofpacket;                                                             // cmd_xbar_demux_008:src10_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src10_valid;                                                                   // cmd_xbar_demux_008:src10_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src10_startofpacket;                                                           // cmd_xbar_demux_008:src10_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src10_data;                                                                    // cmd_xbar_demux_008:src10_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src10_channel;                                                                 // cmd_xbar_demux_008:src10_channel -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src11_endofpacket;                                                             // cmd_xbar_demux_008:src11_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src11_valid;                                                                   // cmd_xbar_demux_008:src11_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src11_startofpacket;                                                           // cmd_xbar_demux_008:src11_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src11_data;                                                                    // cmd_xbar_demux_008:src11_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src11_channel;                                                                 // cmd_xbar_demux_008:src11_channel -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src12_endofpacket;                                                             // cmd_xbar_demux_008:src12_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src12_valid;                                                                   // cmd_xbar_demux_008:src12_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src12_startofpacket;                                                           // cmd_xbar_demux_008:src12_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src12_data;                                                                    // cmd_xbar_demux_008:src12_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src12_channel;                                                                 // cmd_xbar_demux_008:src12_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src13_endofpacket;                                                             // cmd_xbar_demux_008:src13_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src13_valid;                                                                   // cmd_xbar_demux_008:src13_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src13_startofpacket;                                                           // cmd_xbar_demux_008:src13_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src13_data;                                                                    // cmd_xbar_demux_008:src13_data -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src13_channel;                                                                 // cmd_xbar_demux_008:src13_channel -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src14_endofpacket;                                                             // cmd_xbar_demux_008:src14_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src14_valid;                                                                   // cmd_xbar_demux_008:src14_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src14_startofpacket;                                                           // cmd_xbar_demux_008:src14_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src14_data;                                                                    // cmd_xbar_demux_008:src14_data -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src14_channel;                                                                 // cmd_xbar_demux_008:src14_channel -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src15_endofpacket;                                                             // cmd_xbar_demux_008:src15_endofpacket -> ir_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src15_valid;                                                                   // cmd_xbar_demux_008:src15_valid -> ir_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src15_startofpacket;                                                           // cmd_xbar_demux_008:src15_startofpacket -> ir_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src15_data;                                                                    // cmd_xbar_demux_008:src15_data -> ir_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src15_channel;                                                                 // cmd_xbar_demux_008:src15_channel -> ir_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src16_endofpacket;                                                             // cmd_xbar_demux_008:src16_endofpacket -> rs232_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src16_valid;                                                                   // cmd_xbar_demux_008:src16_valid -> rs232_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src16_startofpacket;                                                           // cmd_xbar_demux_008:src16_startofpacket -> rs232_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src16_data;                                                                    // cmd_xbar_demux_008:src16_data -> rs232_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src16_channel;                                                                 // cmd_xbar_demux_008:src16_channel -> rs232_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src17_endofpacket;                                                             // cmd_xbar_demux_008:src17_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src17_valid;                                                                   // cmd_xbar_demux_008:src17_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src17_startofpacket;                                                           // cmd_xbar_demux_008:src17_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_008_src17_data;                                                                    // cmd_xbar_demux_008:src17_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [17:0] cmd_xbar_demux_008_src17_channel;                                                                 // cmd_xbar_demux_008:src17_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                              // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_008:sink0_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                    // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_008:sink0_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                            // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_008:sink0_startofpacket
	wire   [83:0] rsp_xbar_demux_019_src0_data;                                                                     // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_008:sink0_data
	wire   [17:0] rsp_xbar_demux_019_src0_channel;                                                                  // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_008:sink0_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                    // rsp_xbar_mux_008:sink0_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                              // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_008:sink1_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                    // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_008:sink1_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                            // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_008:sink1_startofpacket
	wire   [83:0] rsp_xbar_demux_020_src0_data;                                                                     // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_008:sink1_data
	wire   [17:0] rsp_xbar_demux_020_src0_channel;                                                                  // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_008:sink1_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                    // rsp_xbar_mux_008:sink1_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                              // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_008:sink2_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                    // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_008:sink2_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                            // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_008:sink2_startofpacket
	wire   [83:0] rsp_xbar_demux_021_src0_data;                                                                     // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_008:sink2_data
	wire   [17:0] rsp_xbar_demux_021_src0_channel;                                                                  // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_008:sink2_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                    // rsp_xbar_mux_008:sink2_ready -> rsp_xbar_demux_021:src0_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                              // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_008:sink3_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                    // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_008:sink3_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                            // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_008:sink3_startofpacket
	wire   [83:0] rsp_xbar_demux_022_src0_data;                                                                     // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_008:sink3_data
	wire   [17:0] rsp_xbar_demux_022_src0_channel;                                                                  // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_008:sink3_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                    // rsp_xbar_mux_008:sink3_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                              // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_008:sink4_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                    // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_008:sink4_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                            // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_008:sink4_startofpacket
	wire   [83:0] rsp_xbar_demux_023_src0_data;                                                                     // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_008:sink4_data
	wire   [17:0] rsp_xbar_demux_023_src0_channel;                                                                  // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_008:sink4_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                    // rsp_xbar_mux_008:sink4_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                              // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_008:sink5_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                    // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_008:sink5_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                            // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_008:sink5_startofpacket
	wire   [83:0] rsp_xbar_demux_024_src0_data;                                                                     // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_008:sink5_data
	wire   [17:0] rsp_xbar_demux_024_src0_channel;                                                                  // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_008:sink5_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                    // rsp_xbar_mux_008:sink5_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                              // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_008:sink6_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                    // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_008:sink6_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                            // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_008:sink6_startofpacket
	wire   [83:0] rsp_xbar_demux_025_src0_data;                                                                     // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_008:sink6_data
	wire   [17:0] rsp_xbar_demux_025_src0_channel;                                                                  // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_008:sink6_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                    // rsp_xbar_mux_008:sink6_ready -> rsp_xbar_demux_025:src0_ready
	wire          rsp_xbar_demux_026_src0_endofpacket;                                                              // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_008:sink7_endofpacket
	wire          rsp_xbar_demux_026_src0_valid;                                                                    // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_008:sink7_valid
	wire          rsp_xbar_demux_026_src0_startofpacket;                                                            // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_008:sink7_startofpacket
	wire   [83:0] rsp_xbar_demux_026_src0_data;                                                                     // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_008:sink7_data
	wire   [17:0] rsp_xbar_demux_026_src0_channel;                                                                  // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_008:sink7_channel
	wire          rsp_xbar_demux_026_src0_ready;                                                                    // rsp_xbar_mux_008:sink7_ready -> rsp_xbar_demux_026:src0_ready
	wire          rsp_xbar_demux_027_src0_endofpacket;                                                              // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_008:sink8_endofpacket
	wire          rsp_xbar_demux_027_src0_valid;                                                                    // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_008:sink8_valid
	wire          rsp_xbar_demux_027_src0_startofpacket;                                                            // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_008:sink8_startofpacket
	wire   [83:0] rsp_xbar_demux_027_src0_data;                                                                     // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_008:sink8_data
	wire   [17:0] rsp_xbar_demux_027_src0_channel;                                                                  // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_008:sink8_channel
	wire          rsp_xbar_demux_027_src0_ready;                                                                    // rsp_xbar_mux_008:sink8_ready -> rsp_xbar_demux_027:src0_ready
	wire          rsp_xbar_demux_028_src0_endofpacket;                                                              // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_008:sink9_endofpacket
	wire          rsp_xbar_demux_028_src0_valid;                                                                    // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_008:sink9_valid
	wire          rsp_xbar_demux_028_src0_startofpacket;                                                            // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_008:sink9_startofpacket
	wire   [83:0] rsp_xbar_demux_028_src0_data;                                                                     // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_008:sink9_data
	wire   [17:0] rsp_xbar_demux_028_src0_channel;                                                                  // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_008:sink9_channel
	wire          rsp_xbar_demux_028_src0_ready;                                                                    // rsp_xbar_mux_008:sink9_ready -> rsp_xbar_demux_028:src0_ready
	wire          rsp_xbar_demux_029_src0_endofpacket;                                                              // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_008:sink10_endofpacket
	wire          rsp_xbar_demux_029_src0_valid;                                                                    // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_008:sink10_valid
	wire          rsp_xbar_demux_029_src0_startofpacket;                                                            // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_008:sink10_startofpacket
	wire   [83:0] rsp_xbar_demux_029_src0_data;                                                                     // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_008:sink10_data
	wire   [17:0] rsp_xbar_demux_029_src0_channel;                                                                  // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_008:sink10_channel
	wire          rsp_xbar_demux_029_src0_ready;                                                                    // rsp_xbar_mux_008:sink10_ready -> rsp_xbar_demux_029:src0_ready
	wire          rsp_xbar_demux_030_src0_endofpacket;                                                              // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_008:sink11_endofpacket
	wire          rsp_xbar_demux_030_src0_valid;                                                                    // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_008:sink11_valid
	wire          rsp_xbar_demux_030_src0_startofpacket;                                                            // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_008:sink11_startofpacket
	wire   [83:0] rsp_xbar_demux_030_src0_data;                                                                     // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_008:sink11_data
	wire   [17:0] rsp_xbar_demux_030_src0_channel;                                                                  // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_008:sink11_channel
	wire          rsp_xbar_demux_030_src0_ready;                                                                    // rsp_xbar_mux_008:sink11_ready -> rsp_xbar_demux_030:src0_ready
	wire          rsp_xbar_demux_031_src0_endofpacket;                                                              // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_008:sink12_endofpacket
	wire          rsp_xbar_demux_031_src0_valid;                                                                    // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_008:sink12_valid
	wire          rsp_xbar_demux_031_src0_startofpacket;                                                            // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_008:sink12_startofpacket
	wire   [83:0] rsp_xbar_demux_031_src0_data;                                                                     // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_008:sink12_data
	wire   [17:0] rsp_xbar_demux_031_src0_channel;                                                                  // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_008:sink12_channel
	wire          rsp_xbar_demux_031_src0_ready;                                                                    // rsp_xbar_mux_008:sink12_ready -> rsp_xbar_demux_031:src0_ready
	wire          rsp_xbar_demux_032_src0_endofpacket;                                                              // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_008:sink13_endofpacket
	wire          rsp_xbar_demux_032_src0_valid;                                                                    // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_008:sink13_valid
	wire          rsp_xbar_demux_032_src0_startofpacket;                                                            // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_008:sink13_startofpacket
	wire   [83:0] rsp_xbar_demux_032_src0_data;                                                                     // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_008:sink13_data
	wire   [17:0] rsp_xbar_demux_032_src0_channel;                                                                  // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_008:sink13_channel
	wire          rsp_xbar_demux_032_src0_ready;                                                                    // rsp_xbar_mux_008:sink13_ready -> rsp_xbar_demux_032:src0_ready
	wire          rsp_xbar_demux_033_src0_endofpacket;                                                              // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux_008:sink14_endofpacket
	wire          rsp_xbar_demux_033_src0_valid;                                                                    // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux_008:sink14_valid
	wire          rsp_xbar_demux_033_src0_startofpacket;                                                            // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux_008:sink14_startofpacket
	wire   [83:0] rsp_xbar_demux_033_src0_data;                                                                     // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux_008:sink14_data
	wire   [17:0] rsp_xbar_demux_033_src0_channel;                                                                  // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux_008:sink14_channel
	wire          rsp_xbar_demux_033_src0_ready;                                                                    // rsp_xbar_mux_008:sink14_ready -> rsp_xbar_demux_033:src0_ready
	wire          rsp_xbar_demux_034_src0_endofpacket;                                                              // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux_008:sink15_endofpacket
	wire          rsp_xbar_demux_034_src0_valid;                                                                    // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux_008:sink15_valid
	wire          rsp_xbar_demux_034_src0_startofpacket;                                                            // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux_008:sink15_startofpacket
	wire   [83:0] rsp_xbar_demux_034_src0_data;                                                                     // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux_008:sink15_data
	wire   [17:0] rsp_xbar_demux_034_src0_channel;                                                                  // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux_008:sink15_channel
	wire          rsp_xbar_demux_034_src0_ready;                                                                    // rsp_xbar_mux_008:sink15_ready -> rsp_xbar_demux_034:src0_ready
	wire          rsp_xbar_demux_035_src0_endofpacket;                                                              // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux_008:sink16_endofpacket
	wire          rsp_xbar_demux_035_src0_valid;                                                                    // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux_008:sink16_valid
	wire          rsp_xbar_demux_035_src0_startofpacket;                                                            // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux_008:sink16_startofpacket
	wire   [83:0] rsp_xbar_demux_035_src0_data;                                                                     // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux_008:sink16_data
	wire   [17:0] rsp_xbar_demux_035_src0_channel;                                                                  // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux_008:sink16_channel
	wire          rsp_xbar_demux_035_src0_ready;                                                                    // rsp_xbar_mux_008:sink16_ready -> rsp_xbar_demux_035:src0_ready
	wire          rsp_xbar_demux_036_src0_endofpacket;                                                              // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux_008:sink17_endofpacket
	wire          rsp_xbar_demux_036_src0_valid;                                                                    // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux_008:sink17_valid
	wire          rsp_xbar_demux_036_src0_startofpacket;                                                            // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux_008:sink17_startofpacket
	wire   [83:0] rsp_xbar_demux_036_src0_data;                                                                     // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux_008:sink17_data
	wire   [17:0] rsp_xbar_demux_036_src0_channel;                                                                  // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux_008:sink17_channel
	wire          rsp_xbar_demux_036_src0_ready;                                                                    // rsp_xbar_mux_008:sink17_ready -> rsp_xbar_demux_036:src0_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                  // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire   [83:0] limiter_002_cmd_src_data;                                                                         // limiter_002:cmd_src_data -> cmd_xbar_demux_008:sink_data
	wire   [17:0] limiter_002_cmd_src_channel;                                                                      // limiter_002:cmd_src_channel -> cmd_xbar_demux_008:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                        // cmd_xbar_demux_008:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_008_src_endofpacket;                                                                 // rsp_xbar_mux_008:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_008_src_valid;                                                                       // rsp_xbar_mux_008:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_008_src_startofpacket;                                                               // rsp_xbar_mux_008:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire   [83:0] rsp_xbar_mux_008_src_data;                                                                        // rsp_xbar_mux_008:src_data -> limiter_002:rsp_sink_data
	wire   [17:0] rsp_xbar_mux_008_src_channel;                                                                     // rsp_xbar_mux_008:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_008_src_ready;                                                                       // limiter_002:rsp_sink_ready -> rsp_xbar_mux_008:src_ready
	wire          cmd_xbar_demux_008_src0_ready;                                                                    // key_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src0_ready
	wire          id_router_019_src_endofpacket;                                                                    // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                          // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                  // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire   [83:0] id_router_019_src_data;                                                                           // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [17:0] id_router_019_src_channel;                                                                        // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                          // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_008_src1_ready;                                                                    // lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src1_ready
	wire          id_router_020_src_endofpacket;                                                                    // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                          // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                  // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire   [83:0] id_router_020_src_data;                                                                           // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [17:0] id_router_020_src_channel;                                                                        // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                          // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_008_src2_ready;                                                                    // sd_clk_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src2_ready
	wire          id_router_021_src_endofpacket;                                                                    // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                          // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                  // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire   [83:0] id_router_021_src_data;                                                                           // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [17:0] id_router_021_src_channel;                                                                        // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                          // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          cmd_xbar_demux_008_src3_ready;                                                                    // sd_cmd_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src3_ready
	wire          id_router_022_src_endofpacket;                                                                    // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                          // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                  // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire   [83:0] id_router_022_src_data;                                                                           // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [17:0] id_router_022_src_channel;                                                                        // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                          // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_008_src4_ready;                                                                    // sd_dat_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src4_ready
	wire          id_router_023_src_endofpacket;                                                                    // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                          // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                  // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire   [83:0] id_router_023_src_data;                                                                           // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [17:0] id_router_023_src_channel;                                                                        // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                          // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_demux_008_src5_ready;                                                                    // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src5_ready
	wire          id_router_024_src_endofpacket;                                                                    // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                          // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                  // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire   [83:0] id_router_024_src_data;                                                                           // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [17:0] id_router_024_src_channel;                                                                        // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                          // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_demux_008_src6_ready;                                                                    // epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src6_ready
	wire          id_router_025_src_endofpacket;                                                                    // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                          // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                  // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire   [83:0] id_router_025_src_data;                                                                           // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire   [17:0] id_router_025_src_channel;                                                                        // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                          // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          cmd_xbar_demux_008_src7_ready;                                                                    // epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src7_ready
	wire          id_router_026_src_endofpacket;                                                                    // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire          id_router_026_src_valid;                                                                          // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire          id_router_026_src_startofpacket;                                                                  // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire   [83:0] id_router_026_src_data;                                                                           // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire   [17:0] id_router_026_src_channel;                                                                        // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire          id_router_026_src_ready;                                                                          // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire          cmd_xbar_demux_008_src8_ready;                                                                    // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src8_ready
	wire          id_router_027_src_endofpacket;                                                                    // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire          id_router_027_src_valid;                                                                          // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire          id_router_027_src_startofpacket;                                                                  // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire   [83:0] id_router_027_src_data;                                                                           // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire   [17:0] id_router_027_src_channel;                                                                        // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire          id_router_027_src_ready;                                                                          // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire          cmd_xbar_demux_008_src9_ready;                                                                    // sw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src9_ready
	wire          id_router_028_src_endofpacket;                                                                    // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire          id_router_028_src_valid;                                                                          // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire          id_router_028_src_startofpacket;                                                                  // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire   [83:0] id_router_028_src_data;                                                                           // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire   [17:0] id_router_028_src_channel;                                                                        // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire          id_router_028_src_ready;                                                                          // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire          cmd_xbar_demux_008_src10_ready;                                                                   // i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src10_ready
	wire          id_router_029_src_endofpacket;                                                                    // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire          id_router_029_src_valid;                                                                          // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire          id_router_029_src_startofpacket;                                                                  // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire   [83:0] id_router_029_src_data;                                                                           // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire   [17:0] id_router_029_src_channel;                                                                        // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire          id_router_029_src_ready;                                                                          // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire          cmd_xbar_demux_008_src11_ready;                                                                   // i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src11_ready
	wire          id_router_030_src_endofpacket;                                                                    // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire          id_router_030_src_valid;                                                                          // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire          id_router_030_src_startofpacket;                                                                  // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire   [83:0] id_router_030_src_data;                                                                           // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire   [17:0] id_router_030_src_channel;                                                                        // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire          id_router_030_src_ready;                                                                          // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire          cmd_xbar_demux_008_src12_ready;                                                                   // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src12_ready
	wire          id_router_031_src_endofpacket;                                                                    // id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire          id_router_031_src_valid;                                                                          // id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	wire          id_router_031_src_startofpacket;                                                                  // id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire   [83:0] id_router_031_src_data;                                                                           // id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	wire   [17:0] id_router_031_src_channel;                                                                        // id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	wire          id_router_031_src_ready;                                                                          // rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	wire          cmd_xbar_demux_008_src13_ready;                                                                   // ledg_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src13_ready
	wire          id_router_032_src_endofpacket;                                                                    // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire          id_router_032_src_valid;                                                                          // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire          id_router_032_src_startofpacket;                                                                  // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire   [83:0] id_router_032_src_data;                                                                           // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire   [17:0] id_router_032_src_channel;                                                                        // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire          id_router_032_src_ready;                                                                          // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire          cmd_xbar_demux_008_src14_ready;                                                                   // ledr_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src14_ready
	wire          id_router_033_src_endofpacket;                                                                    // id_router_033:src_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire          id_router_033_src_valid;                                                                          // id_router_033:src_valid -> rsp_xbar_demux_033:sink_valid
	wire          id_router_033_src_startofpacket;                                                                  // id_router_033:src_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire   [83:0] id_router_033_src_data;                                                                           // id_router_033:src_data -> rsp_xbar_demux_033:sink_data
	wire   [17:0] id_router_033_src_channel;                                                                        // id_router_033:src_channel -> rsp_xbar_demux_033:sink_channel
	wire          id_router_033_src_ready;                                                                          // rsp_xbar_demux_033:sink_ready -> id_router_033:src_ready
	wire          cmd_xbar_demux_008_src15_ready;                                                                   // ir_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src15_ready
	wire          id_router_034_src_endofpacket;                                                                    // id_router_034:src_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire          id_router_034_src_valid;                                                                          // id_router_034:src_valid -> rsp_xbar_demux_034:sink_valid
	wire          id_router_034_src_startofpacket;                                                                  // id_router_034:src_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire   [83:0] id_router_034_src_data;                                                                           // id_router_034:src_data -> rsp_xbar_demux_034:sink_data
	wire   [17:0] id_router_034_src_channel;                                                                        // id_router_034:src_channel -> rsp_xbar_demux_034:sink_channel
	wire          id_router_034_src_ready;                                                                          // rsp_xbar_demux_034:sink_ready -> id_router_034:src_ready
	wire          cmd_xbar_demux_008_src16_ready;                                                                   // rs232_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src16_ready
	wire          id_router_035_src_endofpacket;                                                                    // id_router_035:src_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire          id_router_035_src_valid;                                                                          // id_router_035:src_valid -> rsp_xbar_demux_035:sink_valid
	wire          id_router_035_src_startofpacket;                                                                  // id_router_035:src_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire   [83:0] id_router_035_src_data;                                                                           // id_router_035:src_data -> rsp_xbar_demux_035:sink_data
	wire   [17:0] id_router_035_src_channel;                                                                        // id_router_035:src_channel -> rsp_xbar_demux_035:sink_channel
	wire          id_router_035_src_ready;                                                                          // rsp_xbar_demux_035:sink_ready -> id_router_035:src_ready
	wire          cmd_xbar_demux_008_src17_ready;                                                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src17_ready
	wire          id_router_036_src_endofpacket;                                                                    // id_router_036:src_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire          id_router_036_src_valid;                                                                          // id_router_036:src_valid -> rsp_xbar_demux_036:sink_valid
	wire          id_router_036_src_startofpacket;                                                                  // id_router_036:src_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire   [83:0] id_router_036_src_data;                                                                           // id_router_036:src_data -> rsp_xbar_demux_036:sink_data
	wire   [17:0] id_router_036_src_channel;                                                                        // id_router_036:src_channel -> rsp_xbar_demux_036:sink_channel
	wire          id_router_036_src_ready;                                                                          // rsp_xbar_demux_036:sink_ready -> id_router_036:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                 // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                       // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                               // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [106:0] cmd_xbar_mux_001_src_data;                                                                        // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire   [18:0] cmd_xbar_mux_001_src_channel;                                                                     // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire          width_adapter_src_endofpacket;                                                                    // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                          // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                  // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [79:0] width_adapter_src_data;                                                                           // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                          // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [18:0] width_adapter_src_channel;                                                                        // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_001_src_valid;                                                                          // id_router_001:src_valid -> width_adapter_001:in_valid
	wire          id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [79:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> width_adapter_001:in_data
	wire   [18:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> width_adapter_001:in_channel
	wire          id_router_001_src_ready;                                                                          // width_adapter_001:in_ready -> id_router_001:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                      // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                              // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [106:0] width_adapter_001_src_data;                                                                       // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_001_src_ready;                                                                      // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [18:0] width_adapter_001_src_channel;                                                                    // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                 // cmd_xbar_mux_004:src_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                       // cmd_xbar_mux_004:src_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                               // cmd_xbar_mux_004:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [106:0] cmd_xbar_mux_004_src_data;                                                                        // cmd_xbar_mux_004:src_data -> width_adapter_002:in_data
	wire   [18:0] cmd_xbar_mux_004_src_channel;                                                                     // cmd_xbar_mux_004:src_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                       // width_adapter_002:in_ready -> cmd_xbar_mux_004:src_ready
	wire          width_adapter_002_src_endofpacket;                                                                // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                      // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                              // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [88:0] width_adapter_002_src_data;                                                                       // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                      // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire   [18:0] width_adapter_002_src_channel;                                                                    // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_004_src_endofpacket;                                                                    // id_router_004:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_004_src_valid;                                                                          // id_router_004:src_valid -> width_adapter_003:in_valid
	wire          id_router_004_src_startofpacket;                                                                  // id_router_004:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [88:0] id_router_004_src_data;                                                                           // id_router_004:src_data -> width_adapter_003:in_data
	wire   [18:0] id_router_004_src_channel;                                                                        // id_router_004:src_channel -> width_adapter_003:in_channel
	wire          id_router_004_src_ready;                                                                          // width_adapter_003:in_ready -> id_router_004:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                // width_adapter_003:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                      // width_adapter_003:out_valid -> rsp_xbar_demux_004:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                              // width_adapter_003:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] width_adapter_003_src_data;                                                                       // width_adapter_003:out_data -> rsp_xbar_demux_004:sink_data
	wire          width_adapter_003_src_ready;                                                                      // rsp_xbar_demux_004:sink_ready -> width_adapter_003:out_ready
	wire   [18:0] width_adapter_003_src_channel;                                                                    // width_adapter_003:out_channel -> rsp_xbar_demux_004:sink_channel
	wire          crosser_out_endofpacket;                                                                          // crosser:out_endofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                // crosser:out_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                        // crosser:out_startofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] crosser_out_data;                                                                                 // crosser:out_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] crosser_out_channel;                                                                              // crosser:out_channel -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                              // cmd_xbar_demux_001:src8_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                    // cmd_xbar_demux_001:src8_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                            // cmd_xbar_demux_001:src8_startofpacket -> crosser:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src8_data;                                                                     // cmd_xbar_demux_001:src8_data -> crosser:in_data
	wire   [18:0] cmd_xbar_demux_001_src8_channel;                                                                  // cmd_xbar_demux_001:src8_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src8_ready;                                                                    // crosser:in_ready -> cmd_xbar_demux_001:src8_ready
	wire          crosser_001_out_endofpacket;                                                                      // crosser_001:out_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_001_out_valid;                                                                            // crosser_001:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_001_out_startofpacket;                                                                    // crosser_001:out_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] crosser_001_out_data;                                                                             // crosser_001:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] crosser_001_out_channel;                                                                          // crosser_001:out_channel -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                             // cmd_xbar_demux_001:src17_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                   // cmd_xbar_demux_001:src17_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                           // cmd_xbar_demux_001:src17_startofpacket -> crosser_001:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src17_data;                                                                    // cmd_xbar_demux_001:src17_data -> crosser_001:in_data
	wire   [18:0] cmd_xbar_demux_001_src17_channel;                                                                 // cmd_xbar_demux_001:src17_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_001_src17_ready;                                                                   // crosser_001:in_ready -> cmd_xbar_demux_001:src17_ready
	wire          crosser_002_out_endofpacket;                                                                      // crosser_002:out_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_002_out_valid;                                                                            // crosser_002:out_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_002_out_startofpacket;                                                                    // crosser_002:out_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] crosser_002_out_data;                                                                             // crosser_002:out_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] crosser_002_out_channel;                                                                          // crosser_002:out_channel -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                             // cmd_xbar_demux_001:src18_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                   // cmd_xbar_demux_001:src18_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                           // cmd_xbar_demux_001:src18_startofpacket -> crosser_002:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src18_data;                                                                    // cmd_xbar_demux_001:src18_data -> crosser_002:in_data
	wire   [18:0] cmd_xbar_demux_001_src18_channel;                                                                 // cmd_xbar_demux_001:src18_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_001_src18_ready;                                                                   // crosser_002:in_ready -> cmd_xbar_demux_001:src18_ready
	wire          crosser_003_out_endofpacket;                                                                      // crosser_003:out_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          crosser_003_out_valid;                                                                            // crosser_003:out_valid -> rsp_xbar_mux_001:sink8_valid
	wire          crosser_003_out_startofpacket;                                                                    // crosser_003:out_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [106:0] crosser_003_out_data;                                                                             // crosser_003:out_data -> rsp_xbar_mux_001:sink8_data
	wire   [18:0] crosser_003_out_channel;                                                                          // crosser_003:out_channel -> rsp_xbar_mux_001:sink8_channel
	wire          crosser_003_out_ready;                                                                            // rsp_xbar_mux_001:sink8_ready -> crosser_003:out_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                              // rsp_xbar_demux_008:src0_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                    // rsp_xbar_demux_008:src0_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                            // rsp_xbar_demux_008:src0_startofpacket -> crosser_003:in_startofpacket
	wire  [106:0] rsp_xbar_demux_008_src0_data;                                                                     // rsp_xbar_demux_008:src0_data -> crosser_003:in_data
	wire   [18:0] rsp_xbar_demux_008_src0_channel;                                                                  // rsp_xbar_demux_008:src0_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                    // crosser_003:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          crosser_004_out_endofpacket;                                                                      // crosser_004:out_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          crosser_004_out_valid;                                                                            // crosser_004:out_valid -> rsp_xbar_mux_001:sink17_valid
	wire          crosser_004_out_startofpacket;                                                                    // crosser_004:out_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [106:0] crosser_004_out_data;                                                                             // crosser_004:out_data -> rsp_xbar_mux_001:sink17_data
	wire   [18:0] crosser_004_out_channel;                                                                          // crosser_004:out_channel -> rsp_xbar_mux_001:sink17_channel
	wire          crosser_004_out_ready;                                                                            // rsp_xbar_mux_001:sink17_ready -> crosser_004:out_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                              // rsp_xbar_demux_017:src0_endofpacket -> crosser_004:in_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                    // rsp_xbar_demux_017:src0_valid -> crosser_004:in_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                            // rsp_xbar_demux_017:src0_startofpacket -> crosser_004:in_startofpacket
	wire  [106:0] rsp_xbar_demux_017_src0_data;                                                                     // rsp_xbar_demux_017:src0_data -> crosser_004:in_data
	wire   [18:0] rsp_xbar_demux_017_src0_channel;                                                                  // rsp_xbar_demux_017:src0_channel -> crosser_004:in_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                    // crosser_004:in_ready -> rsp_xbar_demux_017:src0_ready
	wire          crosser_005_out_endofpacket;                                                                      // crosser_005:out_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          crosser_005_out_valid;                                                                            // crosser_005:out_valid -> rsp_xbar_mux_001:sink18_valid
	wire          crosser_005_out_startofpacket;                                                                    // crosser_005:out_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [106:0] crosser_005_out_data;                                                                             // crosser_005:out_data -> rsp_xbar_mux_001:sink18_data
	wire   [18:0] crosser_005_out_channel;                                                                          // crosser_005:out_channel -> rsp_xbar_mux_001:sink18_channel
	wire          crosser_005_out_ready;                                                                            // rsp_xbar_mux_001:sink18_ready -> crosser_005:out_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                              // rsp_xbar_demux_018:src0_endofpacket -> crosser_005:in_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                    // rsp_xbar_demux_018:src0_valid -> crosser_005:in_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                            // rsp_xbar_demux_018:src0_startofpacket -> crosser_005:in_startofpacket
	wire  [106:0] rsp_xbar_demux_018_src0_data;                                                                     // rsp_xbar_demux_018:src0_data -> crosser_005:in_data
	wire   [18:0] rsp_xbar_demux_018_src0_channel;                                                                  // rsp_xbar_demux_018:src0_channel -> crosser_005:in_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                    // crosser_005:in_ready -> rsp_xbar_demux_018:src0_ready
	wire   [18:0] limiter_cmd_valid_data;                                                                           // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [18:0] limiter_001_cmd_valid_data;                                                                       // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire   [17:0] limiter_002_cmd_valid_data;                                                                       // limiter_002:cmd_src_valid -> cmd_xbar_demux_008:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                         // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver5_irq;                                                                         // sgdma_tx:csr_irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                                         // sgdma_rx:csr_irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                                                         // ISP1362_IF_0:avs_hc_irq_n_oINT0_N -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                                                         // ISP1362_IF_0:avs_dc_irq_n_oINT0_N -> irq_mapper:receiver8_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                    // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver1_irq;                                                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                    // key:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                         // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                // sw:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver3_irq;                                                                         // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                                // rs232:irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver4_irq;                                                                         // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                                                                // timer:irq -> irq_synchronizer_003:receiver_irq

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (c2_out_clk_clk),                                                    //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                                    // m0_reset.reset
		.s0_clk           (c0_out_clk_clk),                                                    //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (clock_crossing_io_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (clock_crossing_io_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (clock_crossing_io_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (clock_crossing_io_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (clock_crossing_io_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (clock_crossing_io_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (clock_crossing_io_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (clock_crossing_io_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (clock_crossing_io_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (clock_crossing_io_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                                    //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                                      //         .address
		.m0_write         (clock_crossing_io_m0_write),                                        //         .write
		.m0_read          (clock_crossing_io_m0_read),                                         //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                                   //         .debugaccess
	);

	de2_115_WEB_Qsys_cpu cpu (
		.clk                                   (c0_out_clk_clk),                                                     //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	de2_115_WEB_Qsys_tri_state_bridge_flash_bridge_0 tri_state_bridge_flash_bridge_0 (
		.clk                                   (c0_out_clk_clk),                                                           //   clk.clk
		.reset                                 (rst_controller_001_reset_out_reset),                                       // reset.reset
		.request                               (tri_state_flash_bridge_pinsharer_0_tcm_request),                           //   tcs.request
		.grant                                 (tri_state_flash_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.tcs_address_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out),      //      .address_to_the_cfi_flash_out
		.tcs_tri_state_bridge_flash_data       (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out),   //      .tri_state_bridge_flash_data_out
		.tcs_tri_state_bridge_flash_data_outen (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen), //      .tri_state_bridge_flash_data_outen
		.tcs_tri_state_bridge_flash_data_in    (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in),    //      .tri_state_bridge_flash_data_in
		.tcs_write_n_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),      //      .write_n_to_the_cfi_flash_out
		.tcs_select_n_to_the_cfi_flash         (tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),     //      .select_n_to_the_cfi_flash_out
		.tcs_read_n_to_the_cfi_flash           (tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),       //      .read_n_to_the_cfi_flash_out
		.address_to_the_cfi_flash              (tri_state_bridge_flash_bridge_0_out_address_to_the_cfi_flash),             //   out.address_to_the_cfi_flash
		.tri_state_bridge_flash_data           (tri_state_bridge_flash_bridge_0_out_tri_state_bridge_flash_data),          //      .tri_state_bridge_flash_data
		.write_n_to_the_cfi_flash              (tri_state_bridge_flash_bridge_0_out_write_n_to_the_cfi_flash),             //      .write_n_to_the_cfi_flash
		.select_n_to_the_cfi_flash             (tri_state_bridge_flash_bridge_0_out_select_n_to_the_cfi_flash),            //      .select_n_to_the_cfi_flash
		.read_n_to_the_cfi_flash               (tri_state_bridge_flash_bridge_0_out_read_n_to_the_cfi_flash)               //      .read_n_to_the_cfi_flash
	);

	de2_115_WEB_Qsys_tri_state_flash_bridge_pinSharer_0 tri_state_flash_bridge_pinsharer_0 (
		.clk_clk                           (c0_out_clk_clk),                                                           //   clk.clk
		.reset_reset                       (rst_controller_001_reset_out_reset),                                       // reset.reset
		.request                           (tri_state_flash_bridge_pinsharer_0_tcm_request),                           //   tcm.request
		.grant                             (tri_state_flash_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.address_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out),      //      .address_to_the_cfi_flash_out
		.read_n_to_the_cfi_flash           (tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),       //      .read_n_to_the_cfi_flash_out
		.write_n_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),      //      .write_n_to_the_cfi_flash_out
		.tri_state_bridge_flash_data       (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out),   //      .tri_state_bridge_flash_data_out
		.tri_state_bridge_flash_data_in    (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in),    //      .tri_state_bridge_flash_data_in
		.tri_state_bridge_flash_data_outen (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen), //      .tri_state_bridge_flash_data_outen
		.select_n_to_the_cfi_flash         (tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),     //      .select_n_to_the_cfi_flash_out
		.tcs0_request                      (cfi_flash_tcm_request),                                                    //  tcs0.request
		.tcs0_grant                        (cfi_flash_tcm_grant),                                                      //      .grant
		.tcs0_address_out                  (cfi_flash_tcm_address_out),                                                //      .address_out
		.tcs0_read_n_out                   (cfi_flash_tcm_read_n_out),                                                 //      .read_n_out
		.tcs0_write_n_out                  (cfi_flash_tcm_write_n_out),                                                //      .write_n_out
		.tcs0_data_out                     (cfi_flash_tcm_data_out),                                                   //      .data_out
		.tcs0_data_in                      (cfi_flash_tcm_data_in),                                                    //      .data_in
		.tcs0_data_outen                   (cfi_flash_tcm_data_outen),                                                 //      .data_outen
		.tcs0_chipselect_n_out             (cfi_flash_tcm_chipselect_n_out)                                            //      .chipselect_n_out
	);

	de2_115_WEB_Qsys_cfi_flash #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (60),
		.TCM_DATA_HOLD                  (60),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash (
		.clk_clk              (c0_out_clk_clk),                                             //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),                         // reset.reset
		.uas_address          (cfi_flash_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (cfi_flash_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (cfi_flash_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (cfi_flash_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (cfi_flash_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (cfi_flash_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (cfi_flash_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (cfi_flash_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (cfi_flash_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (cfi_flash_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (cfi_flash_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (cfi_flash_tcm_request),                                      //      .request
		.tcm_grant            (cfi_flash_tcm_grant),                                        //      .grant
		.tcm_address_out      (cfi_flash_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (cfi_flash_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (cfi_flash_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (cfi_flash_tcm_data_in)                                       //      .data_in
	);

	de2_115_WEB_Qsys_jtag_uart jtag_uart (
		.clk            (c0_out_clk_clk),                                                         //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	de2_115_WEB_Qsys_key key (
		.clk        (c2_out_clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (key_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~key_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (key_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (key_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (key_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),                   // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)                     //                 irq.irq
	);

	de2_115_WEB_Qsys_lcd lcd (
		.clk           (c2_out_clk_clk),                                                 //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                //         reset.reset_n
		.address       (lcd_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.read          (lcd_control_slave_translator_avalon_anti_slave_0_read),          //              .read
		.readdata      (lcd_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (lcd_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (lcd_control_slave_translator_avalon_anti_slave_0_writedata),     //              .writedata
		.LCD_data      (lcd_external_data),                                              //      external.export
		.LCD_E         (lcd_external_E),                                                 //              .export
		.LCD_RS        (lcd_external_RS),                                                //              .export
		.LCD_RW        (lcd_external_RW)                                                 //              .export
	);

	de2_115_WEB_Qsys_sd_clk sd_clk (
		.clk        (c2_out_clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_clk_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_clk_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_clk_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_clk_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_clk_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (sd_clk_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_sd_cmd sd_cmd (
		.clk        (c2_out_clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_cmd_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_cmd_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_cmd_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_cmd_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_cmd_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (sd_cmd_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_sd_dat sd_dat (
		.clk        (c2_out_clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_dat_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_dat_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_dat_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_dat_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_dat_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (sd_dat_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_sd_wp_n sd_wp_n (
		.clk      (c2_out_clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address  (sd_wp_n_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (sd_wp_n_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (sd_wp_n_external_connection_export)                  // external_connection.export
	);

	de2_115_WEB_Qsys_sd_clk epp_i2c_scl (
		.clk        (c2_out_clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                      //               reset.reset_n
		.address    (epp_i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~epp_i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (epp_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (epp_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (epp_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (epp_i2c_scl_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_sd_cmd epp_i2c_sda (
		.clk        (c2_out_clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (epp_i2c_sda_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~epp_i2c_sda_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (epp_i2c_sda_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (epp_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (epp_i2c_sda_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (epp_i2c_sda_external_connection_export)                    // external_connection.export
	);

	SEG7_IF #(
		.SEG7_NUM       (8),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.s_address   (seg7_avalon_slave_translator_avalon_anti_slave_0_address),   //     avalon_slave.address
		.s_read      (seg7_avalon_slave_translator_avalon_anti_slave_0_read),      //                 .read
		.s_readdata  (seg7_avalon_slave_translator_avalon_anti_slave_0_readdata),  //                 .readdata
		.s_write     (seg7_avalon_slave_translator_avalon_anti_slave_0_write),     //                 .write
		.s_writedata (seg7_avalon_slave_translator_avalon_anti_slave_0_writedata), //                 .writedata
		.SEG7        (seg7_conduit_end_export),                                    //      conduit_end.export
		.s_clk       (c2_out_clk_clk),                                             //       clock_sink.clk
		.s_reset     (rst_controller_reset_out_reset)                              // clock_sink_reset.reset
	);

	de2_115_WEB_Qsys_sw sw (
		.clk        (c2_out_clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (sw_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sw_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sw_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sw_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sw_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),                   // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)                //                 irq.irq
	);

	de2_115_WEB_Qsys_sd_clk i2c_scl (
		.clk        (c2_out_clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_sd_cmd i2c_sda (
		.clk        (c2_out_clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (i2c_sda_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_sda_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)                    // external_connection.export
	);

	AUDIO_IF audio (
		.avs_s1_address       (audio_avalon_slave_translator_avalon_anti_slave_0_address),   //     avalon_slave.address
		.avs_s1_read          (audio_avalon_slave_translator_avalon_anti_slave_0_read),      //                 .read
		.avs_s1_readdata      (audio_avalon_slave_translator_avalon_anti_slave_0_readdata),  //                 .readdata
		.avs_s1_write         (audio_avalon_slave_translator_avalon_anti_slave_0_write),     //                 .write
		.avs_s1_writedata     (audio_avalon_slave_translator_avalon_anti_slave_0_writedata), //                 .writedata
		.avs_s1_clk           (c0_out_clk_clk),                                              //       clock_sink.clk
		.avs_s1_reset         (rst_controller_001_reset_out_reset),                          // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                                       //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                                    //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                                    //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                                    //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                                    //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                                       //                 .export
	);

	de2_115_WEB_Qsys_altpll altpll (
		.clk       (clk_50_clk_in_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_003_reset_out_reset),                        // inclk_interface_reset.reset
		.read      (altpll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (c0_out_clk_clk),                                            //                    c0.clk
		.c1        (altpll_c1_clk),                                             //                    c1.clk
		.c2        (c2_out_clk_clk),                                            //                    c2.clk
		.c3        (altpll_c3_clk),                                             //                    c3.clk
		.areset    (altpll_areset_conduit_export),                              //        areset_conduit.export
		.locked    (altpll_locked_conduit_export),                              //        locked_conduit.export
		.phasedone (altpll_phasedone_conduit_export)                            //     phasedone_conduit.export
	);

	de2_115_WEB_Qsys_onchip_memory2 onchip_memory2 (
		.clk        (c0_out_clk_clk),                                              //   clk1.clk
		.address    (onchip_memory2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                           // reset1.reset
	);

	de2_115_WEB_Qsys_sma_in sma_in (
		.clk      (c0_out_clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address  (sma_in_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (sma_in_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (sma_in_external_connection_export)                  // external_connection.export
	);

	de2_115_WEB_Qsys_sma_out sma_out (
		.clk        (c0_out_clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (sma_out_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sma_out_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sma_out_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sma_out_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sma_out_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (sma_out_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_timer timer (
		.clk        (c2_out_clk_clk),                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_003_receiver_irq)                   //   irq.irq
	);

	de2_115_WEB_Qsys_ledg ledg (
		.clk        (c2_out_clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledg_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledg_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledg_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledg_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledg_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledg_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_ledr ledr (
		.clk        (c2_out_clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)                    // external_connection.export
	);

	de2_115_WEB_Qsys_rs232 rs232 (
		.clk           (c2_out_clk_clk),                                        //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address       (rs232_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (rs232_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (rs232_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~rs232_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~rs232_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (rs232_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (rs232_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                      //                    .dataavailable
		.readyfordata  (),                                                      //                    .readyfordata
		.rxd           (rs232_external_connection_rxd),                         // external_connection.export
		.txd           (rs232_external_connection_txd),                         //                    .export
		.cts_n         (rs232_external_connection_cts_n),                       //                    .export
		.rts_n         (rs232_external_connection_rts_n),                       //                    .export
		.irq           (irq_synchronizer_002_receiver_irq)                      //                 irq.irq
	);

	de2_115_WEB_Qsys_sd_wp_n ir (
		.clk      (c2_out_clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),           //               reset.reset_n
		.address  (ir_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (ir_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (ir_external_connection_export)                  // external_connection.export
	);

	de2_115_WEB_Qsys_sdram sdram (
		.clk            (c0_out_clk_clk),                                        //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	TERASIC_SRAM #(
		.DATA_BITS (16),
		.ADDR_BITS (20)
	) sram (
		.clk            (c0_out_clk_clk),                                               //       clock_reset.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                          // clock_reset_reset.reset_n
		.s_chipselect_n (~sram_avalon_slave_translator_avalon_anti_slave_0_chipselect), //      avalon_slave.chipselect_n
		.s_write_n      (~sram_avalon_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.s_address      (sram_avalon_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.s_read_n       (~sram_avalon_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.s_writedata    (sram_avalon_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.s_readdata     (sram_avalon_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.s_byteenable_n (~sram_avalon_slave_translator_avalon_anti_slave_0_byteenable), //                  .byteenable_n
		.SRAM_DQ        (sram_conduit_end_DQ),                                          //       conduit_end.export
		.SRAM_ADDR      (sram_conduit_end_ADDR),                                        //                  .export
		.SRAM_UB_n      (sram_conduit_end_UB_n),                                        //                  .export
		.SRAM_LB_n      (sram_conduit_end_LB_n),                                        //                  .export
		.SRAM_WE_n      (sram_conduit_end_WE_n),                                        //                  .export
		.SRAM_CE_n      (sram_conduit_end_CE_n),                                        //                  .export
		.SRAM_OE_n      (sram_conduit_end_OE_n)                                         //                  .export
	);

	de2_115_WEB_Qsys_tse_mac tse_mac (
		.ff_tx_data  (sgdma_tx_out_data),                                               //                      transmit.data
		.ff_tx_eop   (sgdma_tx_out_endofpacket),                                        //                              .endofpacket
		.ff_tx_err   (sgdma_tx_out_error),                                              //                              .error
		.ff_tx_mod   (sgdma_tx_out_empty),                                              //                              .empty
		.ff_tx_rdy   (sgdma_tx_out_ready),                                              //                              .ready
		.ff_tx_sop   (sgdma_tx_out_startofpacket),                                      //                              .startofpacket
		.ff_tx_wren  (sgdma_tx_out_valid),                                              //                              .valid
		.ff_tx_clk   (c0_out_clk_clk),                                                  //      receive_clock_connection.clk
		.ff_rx_data  (tse_mac_receive_data),                                            //                       receive.data
		.ff_rx_dval  (tse_mac_receive_valid),                                           //                              .valid
		.ff_rx_eop   (tse_mac_receive_endofpacket),                                     //                              .endofpacket
		.ff_rx_mod   (tse_mac_receive_empty),                                           //                              .empty
		.ff_rx_rdy   (tse_mac_receive_ready),                                           //                              .ready
		.ff_rx_sop   (tse_mac_receive_startofpacket),                                   //                              .startofpacket
		.rx_err      (tse_mac_receive_error),                                           //                              .error
		.ff_rx_clk   (c0_out_clk_clk),                                                  //     transmit_clock_connection.clk
		.address     (tse_mac_control_port_translator_avalon_anti_slave_0_address),     //                  control_port.address
		.readdata    (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),    //                              .readdata
		.read        (tse_mac_control_port_translator_avalon_anti_slave_0_read),        //                              .read
		.writedata   (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),   //                              .writedata
		.write       (tse_mac_control_port_translator_avalon_anti_slave_0_write),       //                              .write
		.waitrequest (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest), //                              .waitrequest
		.clk         (c0_out_clk_clk),                                                  // control_port_clock_connection.clk
		.reset       (rst_controller_001_reset_out_reset),                              //              reset_connection.reset
		.m_rx_d      (tse_mac_conduit_connection_m_rx_d),                               //            conduit_connection.export
		.m_rx_en     (tse_mac_conduit_connection_m_rx_en),                              //                              .export
		.m_rx_err    (tse_mac_conduit_connection_m_rx_err),                             //                              .export
		.m_tx_d      (tse_mac_conduit_connection_m_tx_d),                               //                              .export
		.m_tx_en     (tse_mac_conduit_connection_m_tx_en),                              //                              .export
		.m_tx_err    (tse_mac_conduit_connection_m_tx_err),                             //                              .export
		.tx_clk      (tse_mac_conduit_connection_tx_clk),                               //                              .export
		.rx_clk      (tse_mac_conduit_connection_rx_clk),                               //                              .export
		.set_10      (tse_mac_conduit_connection_set_10),                               //                              .export
		.set_1000    (tse_mac_conduit_connection_set_1000),                             //                              .export
		.ena_10      (tse_mac_conduit_connection_ena_10),                               //                              .export
		.eth_mode    (tse_mac_conduit_connection_eth_mode),                             //                              .export
		.mdio_out    (tse_mac_conduit_connection_mdio_out),                             //                              .export
		.mdio_oen    (tse_mac_conduit_connection_mdio_oen),                             //                              .export
		.mdio_in     (tse_mac_conduit_connection_mdio_in),                              //                              .export
		.mdc         (tse_mac_conduit_connection_mdc),                                  //                              .export
		.m_rx_col    (tse_mac_conduit_connection_m_rx_col),                             //                              .export
		.m_rx_crs    (tse_mac_conduit_connection_m_rx_crs)                              //                              .export
	);

	de2_115_WEB_Qsys_sgdma_tx sgdma_tx (
		.clk                           (c0_out_clk_clk),                                         //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.csr_chipselect                (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_tx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_tx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_tx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver5_irq),                               //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                                //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                                   //                 .read
		.out_data                      (sgdma_tx_out_data),                                      //              out.data
		.out_valid                     (sgdma_tx_out_valid),                                     //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                                     //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                               //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                             //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                                     //                 .empty
		.out_error                     (sgdma_tx_out_error)                                      //                 .error
	);

	de2_115_WEB_Qsys_sgdma_rx sgdma_rx (
		.clk                           (c0_out_clk_clk),                                         //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.csr_chipselect                (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_rx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_rx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_rx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver6_irq),                               //          csr_irq.irq
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),                           //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                               //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                                 //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                             //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable),                            //                 .byteenable
		.in_startofpacket              (tse_mac_receive_startofpacket),                          //               in.startofpacket
		.in_endofpacket                (tse_mac_receive_endofpacket),                            //                 .endofpacket
		.in_empty                      (tse_mac_receive_empty),                                  //                 .empty
		.in_data                       (tse_mac_receive_data),                                   //                 .data
		.in_valid                      (tse_mac_receive_valid),                                  //                 .valid
		.in_ready                      (tse_mac_receive_ready),                                  //                 .ready
		.in_error                      (tse_mac_receive_error)                                   //                 .error
	);

	de2_115_WEB_Qsys_descriptor_memory descriptor_memory (
		.clk        (c0_out_clk_clk),                                                 //   clk1.clk
		.address    (descriptor_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (descriptor_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                              // reset1.reset
	);

	ISP1362_IF isp1362_if_0 (
		.avs_hc_clk_iCLK           (c0_out_clk_clk),                                             //       hc_clock.clk
		.avs_hc_reset_n_iRST_N     (~rst_controller_001_reset_out_reset),                        // hc_clock_reset.reset_n
		.avs_hc_writedata_iDATA    (isp1362_if_0_hc_translator_avalon_anti_slave_0_writedata),   //             hc.writedata
		.avs_hc_readdata_oDATA     (isp1362_if_0_hc_translator_avalon_anti_slave_0_readdata),    //               .readdata
		.avs_hc_address_iADDR      (isp1362_if_0_hc_translator_avalon_anti_slave_0_address),     //               .address
		.avs_hc_read_n_iRD_N       (~isp1362_if_0_hc_translator_avalon_anti_slave_0_read),       //               .read_n
		.avs_hc_write_n_iWR_N      (~isp1362_if_0_hc_translator_avalon_anti_slave_0_write),      //               .write_n
		.avs_hc_chipselect_n_iCS_N (~isp1362_if_0_hc_translator_avalon_anti_slave_0_chipselect), //               .chipselect_n
		.avs_hc_irq_n_oINT0_N      (irq_mapper_receiver7_irq),                                   //         hc_irq.irq_n
		.avs_dc_clk_iCLK           (c0_out_clk_clk),                                             //       dc_clock.clk
		.avs_dc_reset_n_iRST_N     (~cpu_jtag_debug_module_reset_reset),                         // dc_clock_reset.reset_n
		.avs_dc_writedata_iDATA    (isp1362_if_0_dc_translator_avalon_anti_slave_0_writedata),   //             dc.writedata
		.avs_dc_readdata_oDATA     (isp1362_if_0_dc_translator_avalon_anti_slave_0_readdata),    //               .readdata
		.avs_dc_address_iADDR      (isp1362_if_0_dc_translator_avalon_anti_slave_0_address),     //               .address
		.avs_dc_read_n_iRD_N       (~isp1362_if_0_dc_translator_avalon_anti_slave_0_read),       //               .read_n
		.avs_dc_write_n_iWR_N      (~isp1362_if_0_dc_translator_avalon_anti_slave_0_write),      //               .write_n
		.avs_dc_chipselect_n_iCS_N (~isp1362_if_0_dc_translator_avalon_anti_slave_0_chipselect), //               .chipselect_n
		.avs_dc_irq_n_oINT0_N      (irq_mapper_receiver8_irq),                                   //         dc_irq.irq_n
		.USB_DATA                  (isp1362_if_0_conduit_end_DATA),                              //    conduit_end.export
		.USB_ADDR                  (isp1362_if_0_conduit_end_ADDR),                              //               .export
		.USB_RD_N                  (isp1362_if_0_conduit_end_RD_N),                              //               .export
		.USB_WR_N                  (isp1362_if_0_conduit_end_WR_N),                              //               .export
		.USB_CS_N                  (isp1362_if_0_conduit_end_CS_N),                              //               .export
		.USB_RST_N                 (isp1362_if_0_conduit_end_RST_N),                             //               .export
		.USB_INT0                  (isp1362_if_0_conduit_end_INT0),                              //               .export
		.USB_INT1                  (isp1362_if_0_conduit_end_INT1)                               //               .export
	);

	de2_115_WEB_Qsys_sysid sysid (
		.clock    (c2_out_clk_clk),                                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	de2_115_WEB_Qsys_pio_0 pio_0 (
		.clk      (clk_50_clk_in_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_005_reset_out_reset),              //               reset.reset_n
		.address  (pio_0_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_0_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (dataoutput_export)                                 // external_connection.export
	);

	de2_115_WEB_Qsys_pio_1 pio_1 (
		.clk      (clk_50_clk_in_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_005_reset_out_reset),              //               reset.reset_n
		.address  (pio_1_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_1_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (clkoutput_export)                                  // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (c0_out_clk_clk),                                                            //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                        //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (c0_out_clk_clk),                                                     //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_read_translator (
		.clk                   (c0_out_clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_write_translator (
		.clk                   (c0_out_clk_clk),                                                               //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_tx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_tx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_read_translator (
		.clk                   (c0_out_clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_rx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_rx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_rx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_write_translator (
		.clk                   (c0_out_clk_clk),                                                               //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_rx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_m_read_translator (
		.clk                   (c0_out_clk_clk),                                                     //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address           (sgdma_tx_m_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_m_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_m_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_m_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_m_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_m_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_m_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_m_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_write              (1'b0),                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_m_write_translator (
		.clk                   (c0_out_clk_clk),                                                      //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                     reset.reset
		.uav_address           (sgdma_rx_m_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_m_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_m_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_m_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_m_write_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sgdma_rx_m_write_byteenable),                                         //                          .byteenable
		.av_write              (sgdma_rx_m_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_m_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                //               (terminated)
		.av_read               (1'b0),                                                                //               (terminated)
		.av_readdata           (),                                                                    //               (terminated)
		.av_readdatavalid      (),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.av_debugaccess        (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (c0_out_clk_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (23),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cfi_flash_uas_translator (
		.clk                   (c0_out_clk_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cfi_flash_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cfi_flash_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (cfi_flash_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (cfi_flash_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cfi_flash_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (cfi_flash_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (cfi_flash_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (cfi_flash_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (cfi_flash_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (cfi_flash_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (cfi_flash_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_s1_translator (
		.clk                   (c0_out_clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                   (c0_out_clk_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_avalon_slave_translator (
		.clk                   (c0_out_clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_avalon_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (sram_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) clock_crossing_io_s0_translator (
		.clk                   (c0_out_clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (clock_crossing_io_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (clock_crossing_io_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (clock_crossing_io_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (clock_crossing_io_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (clock_crossing_io_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (clock_crossing_io_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (clock_crossing_io_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (clock_crossing_io_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (clock_crossing_io_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (clock_crossing_io_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (c0_out_clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_avalon_slave_translator (
		.clk                   (c0_out_clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_pll_slave_translator (
		.clk                   (clk_50_clk_in_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                          //                    reset.reset
		.uav_address           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (altpll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (altpll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (altpll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (altpll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (altpll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_chipselect         (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sma_in_s1_translator (
		.clk                   (c0_out_clk_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address           (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sma_in_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sma_in_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sma_out_s1_translator (
		.clk                   (c0_out_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sma_out_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sma_out_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sma_out_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sma_out_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sma_out_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (15),
		.AV_WRITE_WAIT_CYCLES           (15),
		.AV_SETUP_WAIT_CYCLES           (15),
		.AV_DATA_HOLD_CYCLES            (15)
	) isp1362_if_0_dc_translator (
		.clk                   (c0_out_clk_clk),                                                             //                      clk.clk
		.reset                 (cpu_jtag_debug_module_reset_reset),                                          //                    reset.reset
		.uav_address           (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (isp1362_if_0_dc_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (isp1362_if_0_dc_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (isp1362_if_0_dc_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (isp1362_if_0_dc_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (isp1362_if_0_dc_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (isp1362_if_0_dc_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_byteenable         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_waitrequest        (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (5),
		.AV_WRITE_WAIT_CYCLES           (5),
		.AV_SETUP_WAIT_CYCLES           (14),
		.AV_DATA_HOLD_CYCLES            (14)
	) isp1362_if_0_hc_translator (
		.clk                   (c0_out_clk_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address           (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (isp1362_if_0_hc_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (isp1362_if_0_hc_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (isp1362_if_0_hc_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (isp1362_if_0_hc_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (isp1362_if_0_hc_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (isp1362_if_0_hc_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_byteenable         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_waitrequest        (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) descriptor_memory_s1_translator (
		.clk                   (c0_out_clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (descriptor_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (descriptor_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_rx_csr_translator (
		.clk                   (c0_out_clk_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_rx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_rx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_rx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_tx_csr_translator (
		.clk                   (c0_out_clk_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_tx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_tx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_tx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tse_mac_control_port_translator (
		.clk                   (c0_out_clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tse_mac_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tse_mac_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (tse_mac_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_0_s1_translator (
		.clk                   (clk_50_clk_in_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                  //                    reset.reset
		.uav_address           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (pio_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                    //              (terminated)
		.av_read               (),                                                                    //              (terminated)
		.av_writedata          (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_chipselect         (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_1_s1_translator (
		.clk                   (clk_50_clk_in_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                  //                    reset.reset
		.uav_address           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (pio_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                    //              (terminated)
		.av_read               (),                                                                    //              (terminated)
		.av_writedata          (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_chipselect         (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (9),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (9),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) clock_crossing_io_m0_translator (
		.clk                   (c2_out_clk_clk),                                                          //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                     reset.reset
		.uav_address           (clock_crossing_io_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (clock_crossing_io_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (clock_crossing_io_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (clock_crossing_io_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (clock_crossing_io_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (clock_crossing_io_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (clock_crossing_io_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (clock_crossing_io_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (clock_crossing_io_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (clock_crossing_io_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (clock_crossing_io_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (clock_crossing_io_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (clock_crossing_io_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (clock_crossing_io_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (clock_crossing_io_m0_byteenable),                                         //                          .byteenable
		.av_read               (clock_crossing_io_m0_read),                                               //                          .read
		.av_readdata           (clock_crossing_io_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (clock_crossing_io_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (clock_crossing_io_m0_write),                                              //                          .write
		.av_writedata          (clock_crossing_io_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (clock_crossing_io_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                    //               (terminated)
		.av_begintransfer      (1'b0),                                                                    //               (terminated)
		.av_chipselect         (1'b0),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                    //               (terminated)
		.uav_clken             (),                                                                        //               (terminated)
		.av_clken              (1'b1)                                                                     //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key_s1_translator (
		.clk                   (c2_out_clk_clk),                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address           (key_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (key_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (key_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (key_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (key_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (key_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (key_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (key_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                  //              (terminated)
		.av_begintransfer      (),                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                  //              (terminated)
		.av_burstcount         (),                                                                  //              (terminated)
		.av_byteenable         (),                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                              //              (terminated)
		.av_writebyteenable    (),                                                                  //              (terminated)
		.av_lock               (),                                                                  //              (terminated)
		.av_clken              (),                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                              //              (terminated)
		.av_debugaccess        (),                                                                  //              (terminated)
		.av_outputenable       ()                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (3),
		.AV_WRITE_WAIT_CYCLES           (3),
		.AV_SETUP_WAIT_CYCLES           (3),
		.AV_DATA_HOLD_CYCLES            (3)
	) lcd_control_slave_translator (
		.clk                   (c2_out_clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lcd_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lcd_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (lcd_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (lcd_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lcd_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_clk_s1_translator (
		.clk                   (c2_out_clk_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_clk_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_clk_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_clk_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_clk_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_clk_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_cmd_s1_translator (
		.clk                   (c2_out_clk_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_cmd_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_cmd_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_cmd_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_cmd_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_cmd_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_dat_s1_translator (
		.clk                   (c2_out_clk_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_dat_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_dat_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_dat_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_dat_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_dat_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_wp_n_s1_translator (
		.clk                   (c2_out_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_wp_n_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sd_wp_n_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                      //              (terminated)
		.av_read               (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epp_i2c_scl_s1_translator (
		.clk                   (c2_out_clk_clk),                                                            //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                        //                    reset.reset
		.uav_address           (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (epp_i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (epp_i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (epp_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (epp_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (epp_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_byteenable         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epp_i2c_sda_s1_translator (
		.clk                   (c2_out_clk_clk),                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address           (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (epp_i2c_sda_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (epp_i2c_sda_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (epp_i2c_sda_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (epp_i2c_sda_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (epp_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_byteenable         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seg7_avalon_slave_translator (
		.clk                   (c2_out_clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (seg7_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (seg7_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (seg7_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (seg7_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (seg7_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sw_s1_translator (
		.clk                   (c2_out_clk_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                   //                    reset.reset
		.uav_address           (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sw_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sw_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sw_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sw_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sw_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                 //              (terminated)
		.av_begintransfer      (),                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                 //              (terminated)
		.av_burstcount         (),                                                                 //              (terminated)
		.av_byteenable         (),                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                             //              (terminated)
		.av_writebyteenable    (),                                                                 //              (terminated)
		.av_lock               (),                                                                 //              (terminated)
		.av_clken              (),                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                             //              (terminated)
		.av_debugaccess        (),                                                                 //              (terminated)
		.av_outputenable       ()                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_scl_s1_translator (
		.clk                   (c2_out_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_sda_s1_translator (
		.clk                   (c2_out_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_sda_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_sda_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                   (c2_out_clk_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledg_s1_translator (
		.clk                   (c2_out_clk_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ledg_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ledg_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ledg_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ledg_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ledg_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledr_s1_translator (
		.clk                   (c2_out_clk_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ir_s1_translator (
		.clk                   (c2_out_clk_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                               //                    reset.reset
		.uav_address           (ir_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ir_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ir_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ir_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ir_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ir_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ir_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (ir_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                 //              (terminated)
		.av_read               (),                                                                 //              (terminated)
		.av_writedata          (),                                                                 //              (terminated)
		.av_begintransfer      (),                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                 //              (terminated)
		.av_burstcount         (),                                                                 //              (terminated)
		.av_byteenable         (),                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                             //              (terminated)
		.av_writebyteenable    (),                                                                 //              (terminated)
		.av_lock               (),                                                                 //              (terminated)
		.av_chipselect         (),                                                                 //              (terminated)
		.av_clken              (),                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                             //              (terminated)
		.av_debugaccess        (),                                                                 //              (terminated)
		.av_outputenable       ()                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rs232_s1_translator (
		.clk                   (c2_out_clk_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (rs232_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rs232_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rs232_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rs232_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rs232_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rs232_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rs232_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rs232_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rs232_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (rs232_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (rs232_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (rs232_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rs232_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rs232_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (rs232_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect         (rs232_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (c2_out_clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                                     //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                              //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                   //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                    //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                 //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src1_valid),                                                        //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src1_data),                                                         //          .data
		.rp_channel       (rsp_xbar_demux_013_src1_channel),                                                      //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src1_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),                                                  //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src1_ready)                                                         //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                                        //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src2_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src2_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_013_src2_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src2_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src2_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src2_ready)                                                          //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src3_valid),                                                        //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src3_data),                                                         //          .data
		.rp_channel       (rsp_xbar_demux_013_src3_channel),                                                      //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src3_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src3_endofpacket),                                                  //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src3_ready)                                                         //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                                        //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src4_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src4_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_013_src4_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src4_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src4_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src4_ready)                                                          //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (6),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_m_read_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                              //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address       (sgdma_tx_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src2_valid),                                               //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src2_data),                                                //          .data
		.rp_channel       (rsp_xbar_demux_003_src2_channel),                                             //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src2_startofpacket),                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),                                         //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src2_ready)                                                //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (7),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_m_write_translator_avalon_universal_master_0_agent (
		.clk              (c0_out_clk_clk),                                                               //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.av_address       (sgdma_rx_m_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_m_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_m_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src3_valid),                                                //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src3_data),                                                 //          .data
		.rp_channel       (rsp_xbar_demux_003_src3_channel),                                              //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src3_startofpacket),                                        //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src3_endofpacket),                                          //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src3_ready)                                                 //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (59),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (60),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (65),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cfi_flash_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                           //                .channel
		.rf_sink_ready           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                  //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (68),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (69),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (74),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                      //                .channel
		.rf_sink_ready           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) clock_crossing_io_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                           //                .channel
		.rf_sink_ready           (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (289),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                         //                .channel
		.rf_sink_ready           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) altpll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_clk_in_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                     //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                     //                .valid
		.cp_data                 (crosser_out_data),                                                                      //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                               //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                   //                .channel
		.rf_sink_ready           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_clk_in_clk),                                                                     //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_50_clk_in_clk),                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.in_data           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sma_in_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sma_in_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                //                .channel
		.rf_sink_ready           (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sma_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sma_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sma_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sma_out_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sma_out_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                //                .channel
		.rf_sink_ready           (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sma_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sma_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sma_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) isp1362_if_0_dc_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                       //             clk.clk
		.reset                   (cpu_jtag_debug_module_reset_reset),                                                    //       clk_reset.reset
		.m0_address              (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                     //                .channel
		.rf_sink_ready           (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                       //       clk.clk
		.reset             (cpu_jtag_debug_module_reset_reset),                                                    // clk_reset.reset
		.in_data           (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) isp1362_if_0_hc_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                     //                .channel
		.rf_sink_ready           (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                              //                .channel
		.rf_sink_ready           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                  //                .channel
		.rf_sink_ready           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                  //                .channel
		.rf_sink_ready           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (c0_out_clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                          //                .channel
		.rf_sink_ready           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c0_out_clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_clk_in_clk),                                                             //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                         //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                         //                .valid
		.cp_data                 (crosser_001_out_data),                                                          //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                   //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                       //                .channel
		.rf_sink_ready           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_clk_in_clk),                                                             //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_50_clk_in_clk),                                                       //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                      // clk_reset.reset
		.in_data           (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_clk_in_clk),                                                             //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                         //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                         //                .valid
		.cp_data                 (crosser_002_out_data),                                                          //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                   //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                       //                .channel
		.rf_sink_ready           (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_clk_in_clk),                                                             //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_50_clk_in_clk),                                                       //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                      // clk_reset.reset
		.in_data           (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.PKT_BURST_TYPE_H          (61),
		.PKT_BURST_TYPE_L          (60),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_TRANS_EXCLUSIVE       (50),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (74),
		.PKT_THREAD_ID_L           (74),
		.PKT_CACHE_H               (81),
		.PKT_CACHE_L               (78),
		.PKT_ADDR_SIDEBAND_H       (62),
		.PKT_ADDR_SIDEBAND_L       (62),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (18),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) clock_crossing_io_m0_translator_avalon_universal_master_0_agent (
		.clk              (c2_out_clk_clk),                                                                   //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (clock_crossing_io_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (clock_crossing_io_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (clock_crossing_io_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (clock_crossing_io_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (clock_crossing_io_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (clock_crossing_io_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (clock_crossing_io_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (clock_crossing_io_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (clock_crossing_io_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (clock_crossing_io_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (clock_crossing_io_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                        //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                         //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                      //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                  //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                         //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) key_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src0_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src0_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_008_src0_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src0_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src0_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src0_channel),                                             //                .channel
		.rf_sink_ready           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src1_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src1_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_008_src1_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src1_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src1_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src1_channel),                                                        //                .channel
		.rf_sink_ready           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_clk_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src2_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src2_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src2_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src2_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src2_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src2_channel),                                                //                .channel
		.rf_sink_ready           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_cmd_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src3_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src3_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src3_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src3_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src3_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src3_channel),                                                //                .channel
		.rf_sink_ready           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_dat_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src4_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src4_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src4_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src4_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src4_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src4_channel),                                                //                .channel
		.rf_sink_ready           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_wp_n_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src5_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src5_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_008_src5_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src5_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src5_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src5_channel),                                                 //                .channel
		.rf_sink_ready           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src6_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src6_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_008_src6_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src6_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src6_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src6_channel),                                                     //                .channel
		.rf_sink_ready           (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src7_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src7_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_008_src7_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src7_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src7_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src7_channel),                                                     //                .channel
		.rf_sink_ready           (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seg7_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src8_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src8_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_008_src8_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src8_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src8_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src8_channel),                                                        //                .channel
		.rf_sink_ready           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sw_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src9_ready),                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src9_valid),                                              //                .valid
		.cp_data                 (cmd_xbar_demux_008_src9_data),                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src9_startofpacket),                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src9_endofpacket),                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src9_channel),                                            //                .channel
		.rf_sink_ready           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.in_data           (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src10_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src10_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src10_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src10_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src10_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src10_channel),                                                //                .channel
		.rf_sink_ready           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src11_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src11_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src11_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src11_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src11_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src11_channel),                                                //                .channel
		.rf_sink_ready           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src12_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src12_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_008_src12_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src12_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src12_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src12_channel),                                              //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ledg_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src13_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src13_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_008_src13_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src13_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src13_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src13_channel),                                             //                .channel
		.rf_sink_ready           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src14_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src14_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_008_src14_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src14_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src14_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src14_channel),                                             //                .channel
		.rf_sink_ready           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ir_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                             //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                         //       clk_reset.reset
		.m0_address              (ir_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ir_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ir_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ir_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ir_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ir_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ir_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ir_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ir_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src15_ready),                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src15_valid),                                             //                .valid
		.cp_data                 (cmd_xbar_demux_008_src15_data),                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src15_startofpacket),                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src15_endofpacket),                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src15_channel),                                           //                .channel
		.rf_sink_ready           (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                             //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                         // clk_reset.reset
		.in_data           (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rs232_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (rs232_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rs232_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rs232_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rs232_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rs232_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rs232_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rs232_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rs232_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rs232_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rs232_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rs232_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rs232_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rs232_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rs232_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src16_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src16_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_008_src16_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src16_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src16_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src16_channel),                                              //                .channel
		.rf_sink_ready           (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (c2_out_clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src17_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src17_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_008_src17_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src17_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src17_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src17_channel),                                                         //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (c2_out_clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	de2_115_WEB_Qsys_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_002 addr_router_002 (
		.sink_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                            //          .valid
		.src_data           (addr_router_002_src_data),                                                             //          .data
		.src_channel        (addr_router_002_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                       //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_002 addr_router_003 (
		.sink_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                             //          .valid
		.src_data           (addr_router_003_src_data),                                                              //          .data
		.src_channel        (addr_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_002 addr_router_004 (
		.sink_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                            //          .valid
		.src_data           (addr_router_004_src_data),                                                             //          .data
		.src_channel        (addr_router_004_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                       //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_002 addr_router_005 (
		.sink_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                             //          .valid
		.src_data           (addr_router_005_src_data),                                                              //          .data
		.src_channel        (addr_router_005_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                        //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_006 addr_router_006 (
		.sink_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                   //          .valid
		.src_data           (addr_router_006_src_data),                                                    //          .data
		.src_channel        (addr_router_006_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                              //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_006 addr_router_007 (
		.sink_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                    //          .valid
		.src_data           (addr_router_007_src_data),                                                     //          .data
		.src_channel        (addr_router_007_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                               //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_001 id_router_001 (
		.sink_ready         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                             //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router id_router_002 (
		.sink_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                      //       src.ready
		.src_valid          (id_router_002_src_valid),                                                      //          .valid
		.src_data           (id_router_002_src_data),                                                       //          .data
		.src_channel        (id_router_002_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                 //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_003 id_router_003 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                             //          .valid
		.src_data           (id_router_003_src_data),                                              //          .data
		.src_channel        (id_router_003_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                        //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_004 id_router_004 (
		.sink_ready         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                      //       src.ready
		.src_valid          (id_router_004_src_valid),                                                      //          .valid
		.src_data           (id_router_004_src_data),                                                       //          .data
		.src_channel        (id_router_004_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                 //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_005 (
		.sink_ready         (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (clock_crossing_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                         //       src.ready
		.src_valid          (id_router_005_src_valid),                                                         //          .valid
		.src_data           (id_router_005_src_data),                                                          //          .data
		.src_channel        (id_router_005_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                    //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_006 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                //          .valid
		.src_data           (id_router_006_src_data),                                                                 //          .data
		.src_channel        (id_router_006_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                           //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_007 (
		.sink_ready         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                       //       src.ready
		.src_valid          (id_router_007_src_valid),                                                       //          .valid
		.src_data           (id_router_007_src_data),                                                        //          .data
		.src_channel        (id_router_007_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                  //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_008 (
		.sink_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_clk_in_clk),                                                           //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                     //       src.ready
		.src_valid          (id_router_008_src_valid),                                                     //          .valid
		.src_data           (id_router_008_src_data),                                                      //          .data
		.src_channel        (id_router_008_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_009 (
		.sink_ready         (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sma_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                              //       src.ready
		.src_valid          (id_router_009_src_valid),                                              //          .valid
		.src_data           (id_router_009_src_data),                                               //          .data
		.src_channel        (id_router_009_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                         //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_010 (
		.sink_ready         (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sma_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                               //          .valid
		.src_data           (id_router_010_src_data),                                                //          .data
		.src_channel        (id_router_010_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                          //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_011 (
		.sink_ready         (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (isp1362_if_0_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                             //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),                                          // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                    //       src.ready
		.src_valid          (id_router_011_src_valid),                                                    //          .valid
		.src_data           (id_router_011_src_data),                                                     //          .data
		.src_channel        (id_router_011_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                               //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_012 (
		.sink_ready         (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (isp1362_if_0_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                    //       src.ready
		.src_valid          (id_router_012_src_valid),                                                    //          .valid
		.src_data           (id_router_012_src_data),                                                     //          .data
		.src_channel        (id_router_012_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                               //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_013 id_router_013 (
		.sink_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                         //       src.ready
		.src_valid          (id_router_013_src_valid),                                                         //          .valid
		.src_data           (id_router_013_src_data),                                                          //          .data
		.src_channel        (id_router_013_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                    //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_014 (
		.sink_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                 //       src.ready
		.src_valid          (id_router_014_src_valid),                                                 //          .valid
		.src_data           (id_router_014_src_data),                                                  //          .data
		.src_channel        (id_router_014_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                            //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_015 (
		.sink_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                 //       src.ready
		.src_valid          (id_router_015_src_valid),                                                 //          .valid
		.src_data           (id_router_015_src_data),                                                  //          .data
		.src_channel        (id_router_015_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                            //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_016 (
		.sink_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c0_out_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                         //       src.ready
		.src_valid          (id_router_016_src_valid),                                                         //          .valid
		.src_data           (id_router_016_src_data),                                                          //          .data
		.src_channel        (id_router_016_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                    //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_017 (
		.sink_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_clk_in_clk),                                                   //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                             //       src.ready
		.src_valid          (id_router_017_src_valid),                                             //          .valid
		.src_data           (id_router_017_src_data),                                              //          .data
		.src_channel        (id_router_017_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                        //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_005 id_router_018 (
		.sink_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_clk_in_clk),                                                   //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                             //       src.ready
		.src_valid          (id_router_018_src_valid),                                             //          .valid
		.src_data           (id_router_018_src_data),                                              //          .data
		.src_channel        (id_router_018_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                        //          .endofpacket
	);

	de2_115_WEB_Qsys_addr_router_008 addr_router_008 (
		.sink_ready         (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (clock_crossing_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                        //          .valid
		.src_data           (addr_router_008_src_data),                                                         //          .data
		.src_channel        (addr_router_008_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                                   //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_019 (
		.sink_ready         (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                           //       src.ready
		.src_valid          (id_router_019_src_valid),                                           //          .valid
		.src_data           (id_router_019_src_data),                                            //          .data
		.src_channel        (id_router_019_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                      //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_020 (
		.sink_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                      //       src.ready
		.src_valid          (id_router_020_src_valid),                                                      //          .valid
		.src_data           (id_router_020_src_data),                                                       //          .data
		.src_channel        (id_router_020_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                 //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_021 (
		.sink_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                              //       src.ready
		.src_valid          (id_router_021_src_valid),                                              //          .valid
		.src_data           (id_router_021_src_data),                                               //          .data
		.src_channel        (id_router_021_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                         //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_022 (
		.sink_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                              //       src.ready
		.src_valid          (id_router_022_src_valid),                                              //          .valid
		.src_data           (id_router_022_src_data),                                               //          .data
		.src_channel        (id_router_022_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                         //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_023 (
		.sink_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                              //       src.ready
		.src_valid          (id_router_023_src_valid),                                              //          .valid
		.src_data           (id_router_023_src_data),                                               //          .data
		.src_channel        (id_router_023_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                         //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_024 (
		.sink_ready         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                               //       src.ready
		.src_valid          (id_router_024_src_valid),                                               //          .valid
		.src_data           (id_router_024_src_data),                                                //          .data
		.src_channel        (id_router_024_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                          //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_025 (
		.sink_ready         (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epp_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                   //       src.ready
		.src_valid          (id_router_025_src_valid),                                                   //          .valid
		.src_data           (id_router_025_src_data),                                                    //          .data
		.src_channel        (id_router_025_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                              //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_026 (
		.sink_ready         (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epp_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                   //       src.ready
		.src_valid          (id_router_026_src_valid),                                                   //          .valid
		.src_data           (id_router_026_src_data),                                                    //          .data
		.src_channel        (id_router_026_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                              //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_027 (
		.sink_ready         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                      //       src.ready
		.src_valid          (id_router_027_src_valid),                                                      //          .valid
		.src_data           (id_router_027_src_data),                                                       //          .data
		.src_channel        (id_router_027_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                                 //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_028 (
		.sink_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                          //       src.ready
		.src_valid          (id_router_028_src_valid),                                          //          .valid
		.src_data           (id_router_028_src_data),                                           //          .data
		.src_channel        (id_router_028_src_channel),                                        //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                     //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_029 (
		.sink_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                               //       src.ready
		.src_valid          (id_router_029_src_valid),                                               //          .valid
		.src_data           (id_router_029_src_data),                                                //          .data
		.src_channel        (id_router_029_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                          //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_030 (
		.sink_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                               //       src.ready
		.src_valid          (id_router_030_src_valid),                                               //          .valid
		.src_data           (id_router_030_src_data),                                                //          .data
		.src_channel        (id_router_030_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                          //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_031 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                             //       src.ready
		.src_valid          (id_router_031_src_valid),                                             //          .valid
		.src_data           (id_router_031_src_data),                                              //          .data
		.src_channel        (id_router_031_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                        //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_032 (
		.sink_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                            //       src.ready
		.src_valid          (id_router_032_src_valid),                                            //          .valid
		.src_data           (id_router_032_src_data),                                             //          .data
		.src_channel        (id_router_032_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                       //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_033 (
		.sink_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                            //       src.ready
		.src_valid          (id_router_033_src_valid),                                            //          .valid
		.src_data           (id_router_033_src_data),                                             //          .data
		.src_channel        (id_router_033_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                       //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_034 (
		.sink_ready         (ir_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ir_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ir_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                               // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                          //       src.ready
		.src_valid          (id_router_034_src_valid),                                          //          .valid
		.src_data           (id_router_034_src_data),                                           //          .data
		.src_channel        (id_router_034_src_channel),                                        //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                     //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_035 (
		.sink_ready         (rs232_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rs232_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rs232_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rs232_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                             //       src.ready
		.src_valid          (id_router_035_src_valid),                                             //          .valid
		.src_data           (id_router_035_src_data),                                              //          .data
		.src_channel        (id_router_035_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                        //          .endofpacket
	);

	de2_115_WEB_Qsys_id_router_019 id_router_036 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (c2_out_clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                                        //       src.ready
		.src_valid          (id_router_036_src_valid),                                                        //          .valid
		.src_data           (id_router_036_src_data),                                                         //          .data
		.src_channel        (id_router_036_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                                   //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (c0_out_clk_clk),                     //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (288),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (c0_out_clk_clk),                     //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (18),
		.VALID_WIDTH               (18),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (c2_out_clk_clk),                     //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_008_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_008_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_008_src_data),           //          .data
		.cmd_sink_channel       (addr_router_008_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_008_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_008_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_008_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_008_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_008_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_008_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_008_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_008_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (59),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (c0_out_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (68),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (c0_out_clk_clk),                          //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (cpu_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                    // reset_in1.reset
		.clk        (c2_out_clk_clk),                    //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.reset_in1  (~reset_reset_n),                     // reset_in1.reset
		.clk        (c0_out_clk_clk),                     //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.clk        (c2_out_clk_clk),                     //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.reset_in1  (~reset_reset_n),                     // reset_in1.reset
		.clk        (clk_50_clk_in_clk),                  //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (c2_out_clk_clk),                     //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_50_clk_in_clk),                  //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	de2_115_WEB_Qsys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (c0_out_clk_clk),                     //        clk.clk
		.reset              (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket)     //           .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (c0_out_clk_clk),                         //        clk.clk
		.reset               (rst_controller_001_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket)    //           .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 cmd_xbar_demux_004 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 cmd_xbar_demux_005 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 cmd_xbar_demux_006 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_006_src_ready),             //      sink.ready
		.sink_channel       (addr_router_006_src_channel),           //          .channel
		.sink_data          (addr_router_006_src_data),              //          .data
		.sink_startofpacket (addr_router_006_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_006_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_006_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 cmd_xbar_demux_007 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_007_src_ready),             //      sink.ready
		.sink_channel       (addr_router_007_src_channel),           //          .channel
		.sink_data          (addr_router_007_src_data),              //          .data
		.sink_startofpacket (addr_router_007_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_007_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_007_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (c0_out_clk_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (c0_out_clk_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (c0_out_clk_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_mux_003 cmd_xbar_mux_003 (
		.clk                 (c0_out_clk_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_006_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_007_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (c0_out_clk_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_mux_013 cmd_xbar_mux_013 (
		.clk                 (c0_out_clk_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src13_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src0_ready),          //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src0_valid),          //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src0_channel),        //          .channel
		.sink3_data          (cmd_xbar_demux_004_src0_data),           //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src0_startofpacket),  //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),    //          .endofpacket
		.sink4_ready         (cmd_xbar_demux_005_src0_ready),          //     sink4.ready
		.sink4_valid         (cmd_xbar_demux_005_src0_valid),          //          .valid
		.sink4_channel       (cmd_xbar_demux_005_src0_channel),        //          .channel
		.sink4_data          (cmd_xbar_demux_005_src0_data),           //          .data
		.sink4_startofpacket (cmd_xbar_demux_005_src0_startofpacket),  //          .startofpacket
		.sink4_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)     //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux rsp_xbar_demux (
		.clk                (c0_out_clk_clk),                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_003_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_003_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_003_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_003_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_003_src3_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (clk_50_clk_in_clk),                     //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),     // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_013 rsp_xbar_demux_013 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_013_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_013_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_013_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_013_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_013_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_013_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_013_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_013_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_013_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_013_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_013_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_013_src3_endofpacket),   //          .endofpacket
		.src4_ready         (rsp_xbar_demux_013_src4_ready),         //      src4.ready
		.src4_valid         (rsp_xbar_demux_013_src4_valid),         //          .valid
		.src4_data          (rsp_xbar_demux_013_src4_data),          //          .data
		.src4_channel       (rsp_xbar_demux_013_src4_channel),       //          .channel
		.src4_startofpacket (rsp_xbar_demux_013_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_013_src4_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_014 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_015 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (c0_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_017 (
		.clk                (clk_50_clk_in_clk),                     //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_002 rsp_xbar_demux_018 (
		.clk                (clk_50_clk_in_clk),                     //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (c0_out_clk_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (c0_out_clk_clk),                        //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (crosser_003_out_ready),                 //     sink8.ready
		.sink8_valid          (crosser_003_out_valid),                 //          .valid
		.sink8_channel        (crosser_003_out_channel),               //          .channel
		.sink8_data           (crosser_003_out_data),                  //          .data
		.sink8_startofpacket  (crosser_003_out_startofpacket),         //          .startofpacket
		.sink8_endofpacket    (crosser_003_out_endofpacket),           //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (crosser_004_out_ready),                 //    sink17.ready
		.sink17_valid         (crosser_004_out_valid),                 //          .valid
		.sink17_channel       (crosser_004_out_channel),               //          .channel
		.sink17_data          (crosser_004_out_data),                  //          .data
		.sink17_startofpacket (crosser_004_out_startofpacket),         //          .startofpacket
		.sink17_endofpacket   (crosser_004_out_endofpacket),           //          .endofpacket
		.sink18_ready         (crosser_005_out_ready),                 //    sink18.ready
		.sink18_valid         (crosser_005_out_valid),                 //          .valid
		.sink18_channel       (crosser_005_out_channel),               //          .channel
		.sink18_data          (crosser_005_out_data),                  //          .data
		.sink18_startofpacket (crosser_005_out_startofpacket),         //          .startofpacket
		.sink18_endofpacket   (crosser_005_out_endofpacket)            //          .endofpacket
	);

	de2_115_WEB_Qsys_cmd_xbar_demux_008 cmd_xbar_demux_008 (
		.clk                 (c2_out_clk_clk),                         //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_002_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_002_cmd_src_channel),            //           .channel
		.sink_data           (limiter_002_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_002_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_002_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_002_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_008_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_008_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_008_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_008_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_008_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_008_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_008_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_008_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_008_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_008_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_008_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_008_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_008_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_008_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_008_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_008_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_008_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_008_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_008_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_008_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_008_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_008_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_008_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_008_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_008_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_008_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_008_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_008_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_008_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_008_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_008_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_008_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_008_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_008_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_008_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_008_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_008_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_008_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_008_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_008_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_008_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_008_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_008_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_008_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_008_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_008_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_008_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_008_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_008_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_008_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_008_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_008_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_008_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_008_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_008_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_008_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_008_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_008_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_008_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_008_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_008_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_008_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_008_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_008_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_008_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_008_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_008_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_008_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_008_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_008_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_008_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_008_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_008_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_008_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_008_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_008_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_008_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_008_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_008_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_008_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_008_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_008_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_008_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_008_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_008_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_008_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_008_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_008_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_008_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_008_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_008_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_008_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_008_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_008_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_008_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_008_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_008_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_008_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_008_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_008_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_008_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_008_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_008_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_008_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_008_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_008_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_008_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_008_src17_endofpacket)    //           .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_019 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_020 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_021 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_022 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_023 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_024 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_025 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_026 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_027 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_028 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_029 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_030 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_031 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_031_src_ready),               //      sink.ready
		.sink_channel       (id_router_031_src_channel),             //          .channel
		.sink_data          (id_router_031_src_data),                //          .data
		.sink_startofpacket (id_router_031_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_031_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_031_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_032 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_033 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_033_src_ready),               //      sink.ready
		.sink_channel       (id_router_033_src_channel),             //          .channel
		.sink_data          (id_router_033_src_data),                //          .data
		.sink_startofpacket (id_router_033_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_033_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_033_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_034 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_034_src_ready),               //      sink.ready
		.sink_channel       (id_router_034_src_channel),             //          .channel
		.sink_data          (id_router_034_src_data),                //          .data
		.sink_startofpacket (id_router_034_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_034_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_034_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_035 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_035_src_ready),               //      sink.ready
		.sink_channel       (id_router_035_src_channel),             //          .channel
		.sink_data          (id_router_035_src_data),                //          .data
		.sink_startofpacket (id_router_035_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_035_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_035_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_demux_019 rsp_xbar_demux_036 (
		.clk                (c2_out_clk_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_036_src_ready),               //      sink.ready
		.sink_channel       (id_router_036_src_channel),             //          .channel
		.sink_data          (id_router_036_src_data),                //          .data
		.sink_startofpacket (id_router_036_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_036_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_036_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	de2_115_WEB_Qsys_rsp_xbar_mux_008 rsp_xbar_mux_008 (
		.clk                  (c2_out_clk_clk),                        //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_008_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_008_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_008_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_019_src0_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_019_src0_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_020_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_020_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_021_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_021_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_022_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_022_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_023_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_023_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_024_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_024_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_025_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_025_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_026_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_026_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_027_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_027_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_028_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_028_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_029_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_030_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_031_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_032_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_033_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_034_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_035_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_036_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (c0_out_clk_clk),                     //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (c0_out_clk_clk),                      //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (c0_out_clk_clk),                      //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (cmd_xbar_mux_004_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_004_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_004_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_004_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_004_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_004_src_data),           //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk                  (c0_out_clk_clk),                      //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_004_src_valid),             //      sink.valid
		.in_channel           (id_router_004_src_channel),           //          .channel
		.in_startofpacket     (id_router_004_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_004_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_004_src_ready),             //          .ready
		.in_data              (id_router_004_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (c0_out_clk_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_50_clk_in_clk),                     //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src8_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src8_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src8_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src8_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src8_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (c0_out_clk_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (clk_50_clk_in_clk),                      //       out_clk.clk
		.out_reset         (rst_controller_005_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src17_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src17_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src17_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src17_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src17_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src17_data),          //              .data
		.out_ready         (crosser_001_out_ready),                  //           out.ready
		.out_valid         (crosser_001_out_valid),                  //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_001_out_channel),                //              .channel
		.out_data          (crosser_001_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (c0_out_clk_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (clk_50_clk_in_clk),                      //       out_clk.clk
		.out_reset         (rst_controller_005_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src18_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src18_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src18_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src18_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src18_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src18_data),          //              .data
		.out_ready         (crosser_002_out_ready),                  //           out.ready
		.out_valid         (crosser_002_out_valid),                  //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_002_out_channel),                //              .channel
		.out_data          (crosser_002_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk_50_clk_in_clk),                     //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (c0_out_clk_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (clk_50_clk_in_clk),                     //        in_clk.clk
		.in_reset          (rst_controller_005_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (c0_out_clk_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_017_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_017_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_017_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_017_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_017_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_017_src0_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (clk_50_clk_in_clk),                     //        in_clk.clk
		.in_reset          (rst_controller_005_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (c0_out_clk_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_018_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_018_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_018_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_018_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_018_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_018_src0_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	de2_115_WEB_Qsys_irq_mapper irq_mapper (
		.clk           (c0_out_clk_clk),                     //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (~irq_mapper_receiver7_irq),          // receiver7.irq
		.receiver8_irq (~irq_mapper_receiver8_irq),          // receiver8.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (c2_out_clk_clk),                     //       receiver_clk.clk
		.sender_clk     (c0_out_clk_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (c2_out_clk_clk),                     //       receiver_clk.clk
		.sender_clk     (c0_out_clk_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (c2_out_clk_clk),                     //       receiver_clk.clk
		.sender_clk     (c0_out_clk_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (c2_out_clk_clk),                     //       receiver_clk.clk
		.sender_clk     (c0_out_clk_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

endmodule
